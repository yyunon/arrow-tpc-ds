-- Copyright 2018-2019 Delft University of Technology
--
-- Licensed under the Apache License, Version 2.0 (the "License");
-- you may not use this file except in compliance with the License.
-- You may obtain a copy of the License at
--
--     http://www.apache.org/licenses/LICENSE-2.0
--
-- Unless required by applicable law or agreed to in writing, software
-- distributed under the License is distributed on an "AS IS" BASIS,
-- WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
-- See the License for the specific language governing permissions and
-- limitations under the License.
--
-- This file was generated by Fletchgen. Modify this file at your own risk.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library work;
use work.Array_pkg.all;

entity Join_ss is
  generic (
    INDEX_WIDTH                        : integer := 32;
    TAG_WIDTH                          : integer := 1;
    SS_SOLD_DATE_SK_BUS_ADDR_WIDTH     : integer := 64;
    SS_SOLD_DATE_SK_BUS_DATA_WIDTH     : integer := 512;
    SS_SOLD_DATE_SK_BUS_LEN_WIDTH      : integer := 8;
    SS_SOLD_DATE_SK_BUS_BURST_STEP_LEN : integer := 1;
    SS_SOLD_DATE_SK_BUS_BURST_MAX_LEN  : integer := 16;
    SS_CDEMO_SK_BUS_ADDR_WIDTH         : integer := 64;
    SS_CDEMO_SK_BUS_DATA_WIDTH         : integer := 512;
    SS_CDEMO_SK_BUS_LEN_WIDTH          : integer := 8;
    SS_CDEMO_SK_BUS_BURST_STEP_LEN     : integer := 1;
    SS_CDEMO_SK_BUS_BURST_MAX_LEN      : integer := 16;
    SS_ADDR_SK_BUS_ADDR_WIDTH          : integer := 64;
    SS_ADDR_SK_BUS_DATA_WIDTH          : integer := 512;
    SS_ADDR_SK_BUS_LEN_WIDTH           : integer := 8;
    SS_ADDR_SK_BUS_BURST_STEP_LEN      : integer := 1;
    SS_ADDR_SK_BUS_BURST_MAX_LEN       : integer := 16;
    SS_STORE_SK_BUS_ADDR_WIDTH         : integer := 64;
    SS_STORE_SK_BUS_DATA_WIDTH         : integer := 512;
    SS_STORE_SK_BUS_LEN_WIDTH          : integer := 8;
    SS_STORE_SK_BUS_BURST_STEP_LEN     : integer := 1;
    SS_STORE_SK_BUS_BURST_MAX_LEN      : integer := 16;
    SS_QUANTITY_BUS_ADDR_WIDTH         : integer := 64;
    SS_QUANTITY_BUS_DATA_WIDTH         : integer := 512;
    SS_QUANTITY_BUS_LEN_WIDTH          : integer := 8;
    SS_QUANTITY_BUS_BURST_STEP_LEN     : integer := 1;
    SS_QUANTITY_BUS_BURST_MAX_LEN      : integer := 16;
    SS_SALES_PRICE_BUS_ADDR_WIDTH      : integer := 64;
    SS_SALES_PRICE_BUS_DATA_WIDTH      : integer := 512;
    SS_SALES_PRICE_BUS_LEN_WIDTH       : integer := 8;
    SS_SALES_PRICE_BUS_BURST_STEP_LEN  : integer := 1;
    SS_SALES_PRICE_BUS_BURST_MAX_LEN   : integer := 16;
    SS_NET_PROFIT_BUS_ADDR_WIDTH       : integer := 64;
    SS_NET_PROFIT_BUS_DATA_WIDTH       : integer := 512;
    SS_NET_PROFIT_BUS_LEN_WIDTH        : integer := 8;
    SS_NET_PROFIT_BUS_BURST_STEP_LEN   : integer := 1;
    SS_NET_PROFIT_BUS_BURST_MAX_LEN    : integer := 16
  );
  port (
    bcd_clk                        : in  std_logic;
    bcd_reset                      : in  std_logic;
    kcd_clk                        : in  std_logic;
    kcd_reset                      : in  std_logic;
    ss_sold_date_sk_valid          : out std_logic;
    ss_sold_date_sk_ready          : in  std_logic;
    ss_sold_date_sk_dvalid         : out std_logic;
    ss_sold_date_sk_last           : out std_logic;
    ss_sold_date_sk                : out std_logic_vector(63 downto 0);
    ss_sold_date_sk_bus_rreq_valid : out std_logic;
    ss_sold_date_sk_bus_rreq_ready : in  std_logic;
    ss_sold_date_sk_bus_rreq_addr  : out std_logic_vector(SS_SOLD_DATE_SK_BUS_ADDR_WIDTH-1 downto 0);
    ss_sold_date_sk_bus_rreq_len   : out std_logic_vector(SS_SOLD_DATE_SK_BUS_LEN_WIDTH-1 downto 0);
    ss_sold_date_sk_bus_rdat_valid : in  std_logic;
    ss_sold_date_sk_bus_rdat_ready : out std_logic;
    ss_sold_date_sk_bus_rdat_data  : in  std_logic_vector(SS_SOLD_DATE_SK_BUS_DATA_WIDTH-1 downto 0);
    ss_sold_date_sk_bus_rdat_last  : in  std_logic;
    ss_sold_date_sk_cmd_valid      : in  std_logic;
    ss_sold_date_sk_cmd_ready      : out std_logic;
    ss_sold_date_sk_cmd_firstIdx   : in  std_logic_vector(INDEX_WIDTH-1 downto 0);
    ss_sold_date_sk_cmd_lastIdx    : in  std_logic_vector(INDEX_WIDTH-1 downto 0);
    ss_sold_date_sk_cmd_ctrl       : in  std_logic_vector(SS_SOLD_DATE_SK_BUS_ADDR_WIDTH-1 downto 0);
    ss_sold_date_sk_cmd_tag        : in  std_logic_vector(TAG_WIDTH-1 downto 0);
    ss_sold_date_sk_unl_valid      : out std_logic;
    ss_sold_date_sk_unl_ready      : in  std_logic;
    ss_sold_date_sk_unl_tag        : out std_logic_vector(TAG_WIDTH-1 downto 0);
    ss_cdemo_sk_valid              : out std_logic;
    ss_cdemo_sk_ready              : in  std_logic;
    ss_cdemo_sk_dvalid             : out std_logic;
    ss_cdemo_sk_last               : out std_logic;
    ss_cdemo_sk                    : out std_logic_vector(63 downto 0);
    ss_cdemo_sk_bus_rreq_valid     : out std_logic;
    ss_cdemo_sk_bus_rreq_ready     : in  std_logic;
    ss_cdemo_sk_bus_rreq_addr      : out std_logic_vector(SS_CDEMO_SK_BUS_ADDR_WIDTH-1 downto 0);
    ss_cdemo_sk_bus_rreq_len       : out std_logic_vector(SS_CDEMO_SK_BUS_LEN_WIDTH-1 downto 0);
    ss_cdemo_sk_bus_rdat_valid     : in  std_logic;
    ss_cdemo_sk_bus_rdat_ready     : out std_logic;
    ss_cdemo_sk_bus_rdat_data      : in  std_logic_vector(SS_CDEMO_SK_BUS_DATA_WIDTH-1 downto 0);
    ss_cdemo_sk_bus_rdat_last      : in  std_logic;
    ss_cdemo_sk_cmd_valid          : in  std_logic;
    ss_cdemo_sk_cmd_ready          : out std_logic;
    ss_cdemo_sk_cmd_firstIdx       : in  std_logic_vector(INDEX_WIDTH-1 downto 0);
    ss_cdemo_sk_cmd_lastIdx        : in  std_logic_vector(INDEX_WIDTH-1 downto 0);
    ss_cdemo_sk_cmd_ctrl           : in  std_logic_vector(SS_CDEMO_SK_BUS_ADDR_WIDTH-1 downto 0);
    ss_cdemo_sk_cmd_tag            : in  std_logic_vector(TAG_WIDTH-1 downto 0);
    ss_cdemo_sk_unl_valid          : out std_logic;
    ss_cdemo_sk_unl_ready          : in  std_logic;
    ss_cdemo_sk_unl_tag            : out std_logic_vector(TAG_WIDTH-1 downto 0);
    ss_addr_sk_valid               : out std_logic;
    ss_addr_sk_ready               : in  std_logic;
    ss_addr_sk_dvalid              : out std_logic;
    ss_addr_sk_last                : out std_logic;
    ss_addr_sk                     : out std_logic_vector(63 downto 0);
    ss_addr_sk_bus_rreq_valid      : out std_logic;
    ss_addr_sk_bus_rreq_ready      : in  std_logic;
    ss_addr_sk_bus_rreq_addr       : out std_logic_vector(SS_ADDR_SK_BUS_ADDR_WIDTH-1 downto 0);
    ss_addr_sk_bus_rreq_len        : out std_logic_vector(SS_ADDR_SK_BUS_LEN_WIDTH-1 downto 0);
    ss_addr_sk_bus_rdat_valid      : in  std_logic;
    ss_addr_sk_bus_rdat_ready      : out std_logic;
    ss_addr_sk_bus_rdat_data       : in  std_logic_vector(SS_ADDR_SK_BUS_DATA_WIDTH-1 downto 0);
    ss_addr_sk_bus_rdat_last       : in  std_logic;
    ss_addr_sk_cmd_valid           : in  std_logic;
    ss_addr_sk_cmd_ready           : out std_logic;
    ss_addr_sk_cmd_firstIdx        : in  std_logic_vector(INDEX_WIDTH-1 downto 0);
    ss_addr_sk_cmd_lastIdx         : in  std_logic_vector(INDEX_WIDTH-1 downto 0);
    ss_addr_sk_cmd_ctrl            : in  std_logic_vector(SS_ADDR_SK_BUS_ADDR_WIDTH-1 downto 0);
    ss_addr_sk_cmd_tag             : in  std_logic_vector(TAG_WIDTH-1 downto 0);
    ss_addr_sk_unl_valid           : out std_logic;
    ss_addr_sk_unl_ready           : in  std_logic;
    ss_addr_sk_unl_tag             : out std_logic_vector(TAG_WIDTH-1 downto 0);
    ss_store_sk_valid              : out std_logic;
    ss_store_sk_ready              : in  std_logic;
    ss_store_sk_dvalid             : out std_logic;
    ss_store_sk_last               : out std_logic;
    ss_store_sk                    : out std_logic_vector(63 downto 0);
    ss_store_sk_bus_rreq_valid     : out std_logic;
    ss_store_sk_bus_rreq_ready     : in  std_logic;
    ss_store_sk_bus_rreq_addr      : out std_logic_vector(SS_STORE_SK_BUS_ADDR_WIDTH-1 downto 0);
    ss_store_sk_bus_rreq_len       : out std_logic_vector(SS_STORE_SK_BUS_LEN_WIDTH-1 downto 0);
    ss_store_sk_bus_rdat_valid     : in  std_logic;
    ss_store_sk_bus_rdat_ready     : out std_logic;
    ss_store_sk_bus_rdat_data      : in  std_logic_vector(SS_STORE_SK_BUS_DATA_WIDTH-1 downto 0);
    ss_store_sk_bus_rdat_last      : in  std_logic;
    ss_store_sk_cmd_valid          : in  std_logic;
    ss_store_sk_cmd_ready          : out std_logic;
    ss_store_sk_cmd_firstIdx       : in  std_logic_vector(INDEX_WIDTH-1 downto 0);
    ss_store_sk_cmd_lastIdx        : in  std_logic_vector(INDEX_WIDTH-1 downto 0);
    ss_store_sk_cmd_ctrl           : in  std_logic_vector(SS_STORE_SK_BUS_ADDR_WIDTH-1 downto 0);
    ss_store_sk_cmd_tag            : in  std_logic_vector(TAG_WIDTH-1 downto 0);
    ss_store_sk_unl_valid          : out std_logic;
    ss_store_sk_unl_ready          : in  std_logic;
    ss_store_sk_unl_tag            : out std_logic_vector(TAG_WIDTH-1 downto 0);
    ss_quantity_valid              : out std_logic;
    ss_quantity_ready              : in  std_logic;
    ss_quantity_dvalid             : out std_logic;
    ss_quantity_last               : out std_logic;
    ss_quantity                    : out std_logic_vector(63 downto 0);
    ss_quantity_bus_rreq_valid     : out std_logic;
    ss_quantity_bus_rreq_ready     : in  std_logic;
    ss_quantity_bus_rreq_addr      : out std_logic_vector(SS_QUANTITY_BUS_ADDR_WIDTH-1 downto 0);
    ss_quantity_bus_rreq_len       : out std_logic_vector(SS_QUANTITY_BUS_LEN_WIDTH-1 downto 0);
    ss_quantity_bus_rdat_valid     : in  std_logic;
    ss_quantity_bus_rdat_ready     : out std_logic;
    ss_quantity_bus_rdat_data      : in  std_logic_vector(SS_QUANTITY_BUS_DATA_WIDTH-1 downto 0);
    ss_quantity_bus_rdat_last      : in  std_logic;
    ss_quantity_cmd_valid          : in  std_logic;
    ss_quantity_cmd_ready          : out std_logic;
    ss_quantity_cmd_firstIdx       : in  std_logic_vector(INDEX_WIDTH-1 downto 0);
    ss_quantity_cmd_lastIdx        : in  std_logic_vector(INDEX_WIDTH-1 downto 0);
    ss_quantity_cmd_ctrl           : in  std_logic_vector(SS_QUANTITY_BUS_ADDR_WIDTH-1 downto 0);
    ss_quantity_cmd_tag            : in  std_logic_vector(TAG_WIDTH-1 downto 0);
    ss_quantity_unl_valid          : out std_logic;
    ss_quantity_unl_ready          : in  std_logic;
    ss_quantity_unl_tag            : out std_logic_vector(TAG_WIDTH-1 downto 0);
    ss_sales_price_valid           : out std_logic;
    ss_sales_price_ready           : in  std_logic;
    ss_sales_price_dvalid          : out std_logic;
    ss_sales_price_last            : out std_logic;
    ss_sales_price                 : out std_logic_vector(63 downto 0);
    ss_sales_price_bus_rreq_valid  : out std_logic;
    ss_sales_price_bus_rreq_ready  : in  std_logic;
    ss_sales_price_bus_rreq_addr   : out std_logic_vector(SS_SALES_PRICE_BUS_ADDR_WIDTH-1 downto 0);
    ss_sales_price_bus_rreq_len    : out std_logic_vector(SS_SALES_PRICE_BUS_LEN_WIDTH-1 downto 0);
    ss_sales_price_bus_rdat_valid  : in  std_logic;
    ss_sales_price_bus_rdat_ready  : out std_logic;
    ss_sales_price_bus_rdat_data   : in  std_logic_vector(SS_SALES_PRICE_BUS_DATA_WIDTH-1 downto 0);
    ss_sales_price_bus_rdat_last   : in  std_logic;
    ss_sales_price_cmd_valid       : in  std_logic;
    ss_sales_price_cmd_ready       : out std_logic;
    ss_sales_price_cmd_firstIdx    : in  std_logic_vector(INDEX_WIDTH-1 downto 0);
    ss_sales_price_cmd_lastIdx     : in  std_logic_vector(INDEX_WIDTH-1 downto 0);
    ss_sales_price_cmd_ctrl        : in  std_logic_vector(SS_SALES_PRICE_BUS_ADDR_WIDTH-1 downto 0);
    ss_sales_price_cmd_tag         : in  std_logic_vector(TAG_WIDTH-1 downto 0);
    ss_sales_price_unl_valid       : out std_logic;
    ss_sales_price_unl_ready       : in  std_logic;
    ss_sales_price_unl_tag         : out std_logic_vector(TAG_WIDTH-1 downto 0);
    ss_net_profit_valid            : out std_logic;
    ss_net_profit_ready            : in  std_logic;
    ss_net_profit_dvalid           : out std_logic;
    ss_net_profit_last             : out std_logic;
    ss_net_profit                  : out std_logic_vector(63 downto 0);
    ss_net_profit_bus_rreq_valid   : out std_logic;
    ss_net_profit_bus_rreq_ready   : in  std_logic;
    ss_net_profit_bus_rreq_addr    : out std_logic_vector(SS_NET_PROFIT_BUS_ADDR_WIDTH-1 downto 0);
    ss_net_profit_bus_rreq_len     : out std_logic_vector(SS_NET_PROFIT_BUS_LEN_WIDTH-1 downto 0);
    ss_net_profit_bus_rdat_valid   : in  std_logic;
    ss_net_profit_bus_rdat_ready   : out std_logic;
    ss_net_profit_bus_rdat_data    : in  std_logic_vector(SS_NET_PROFIT_BUS_DATA_WIDTH-1 downto 0);
    ss_net_profit_bus_rdat_last    : in  std_logic;
    ss_net_profit_cmd_valid        : in  std_logic;
    ss_net_profit_cmd_ready        : out std_logic;
    ss_net_profit_cmd_firstIdx     : in  std_logic_vector(INDEX_WIDTH-1 downto 0);
    ss_net_profit_cmd_lastIdx      : in  std_logic_vector(INDEX_WIDTH-1 downto 0);
    ss_net_profit_cmd_ctrl         : in  std_logic_vector(SS_NET_PROFIT_BUS_ADDR_WIDTH-1 downto 0);
    ss_net_profit_cmd_tag          : in  std_logic_vector(TAG_WIDTH-1 downto 0);
    ss_net_profit_unl_valid        : out std_logic;
    ss_net_profit_unl_ready        : in  std_logic;
    ss_net_profit_unl_tag          : out std_logic_vector(TAG_WIDTH-1 downto 0)
  );
end entity;

architecture Implementation of Join_ss is
  signal sold_date_sk_inst_cmd_valid      : std_logic;
  signal sold_date_sk_inst_cmd_ready      : std_logic;
  signal sold_date_sk_inst_cmd_firstIdx   : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal sold_date_sk_inst_cmd_lastIdx    : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal sold_date_sk_inst_cmd_ctrl       : std_logic_vector(SS_SOLD_DATE_SK_BUS_ADDR_WIDTH-1 downto 0);
  signal sold_date_sk_inst_cmd_tag        : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal sold_date_sk_inst_unl_valid      : std_logic;
  signal sold_date_sk_inst_unl_ready      : std_logic;
  signal sold_date_sk_inst_unl_tag        : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal sold_date_sk_inst_bus_rreq_valid : std_logic;
  signal sold_date_sk_inst_bus_rreq_ready : std_logic;
  signal sold_date_sk_inst_bus_rreq_addr  : std_logic_vector(SS_SOLD_DATE_SK_BUS_ADDR_WIDTH-1 downto 0);
  signal sold_date_sk_inst_bus_rreq_len   : std_logic_vector(SS_SOLD_DATE_SK_BUS_LEN_WIDTH-1 downto 0);
  signal sold_date_sk_inst_bus_rdat_valid : std_logic;
  signal sold_date_sk_inst_bus_rdat_ready : std_logic;
  signal sold_date_sk_inst_bus_rdat_data  : std_logic_vector(SS_SOLD_DATE_SK_BUS_DATA_WIDTH-1 downto 0);
  signal sold_date_sk_inst_bus_rdat_last  : std_logic;

  signal sold_date_sk_inst_out_valid      : std_logic_vector(0 downto 0);
  signal sold_date_sk_inst_out_ready      : std_logic_vector(0 downto 0);
  signal sold_date_sk_inst_out_data       : std_logic_vector(63 downto 0);
  signal sold_date_sk_inst_out_dvalid     : std_logic_vector(0 downto 0);
  signal sold_date_sk_inst_out_last       : std_logic_vector(0 downto 0);

  signal cdemo_sk_inst_cmd_valid          : std_logic;
  signal cdemo_sk_inst_cmd_ready          : std_logic;
  signal cdemo_sk_inst_cmd_firstIdx       : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal cdemo_sk_inst_cmd_lastIdx        : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal cdemo_sk_inst_cmd_ctrl           : std_logic_vector(SS_CDEMO_SK_BUS_ADDR_WIDTH-1 downto 0);
  signal cdemo_sk_inst_cmd_tag            : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal cdemo_sk_inst_unl_valid          : std_logic;
  signal cdemo_sk_inst_unl_ready          : std_logic;
  signal cdemo_sk_inst_unl_tag            : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal cdemo_sk_inst_bus_rreq_valid     : std_logic;
  signal cdemo_sk_inst_bus_rreq_ready     : std_logic;
  signal cdemo_sk_inst_bus_rreq_addr      : std_logic_vector(SS_CDEMO_SK_BUS_ADDR_WIDTH-1 downto 0);
  signal cdemo_sk_inst_bus_rreq_len       : std_logic_vector(SS_CDEMO_SK_BUS_LEN_WIDTH-1 downto 0);
  signal cdemo_sk_inst_bus_rdat_valid     : std_logic;
  signal cdemo_sk_inst_bus_rdat_ready     : std_logic;
  signal cdemo_sk_inst_bus_rdat_data      : std_logic_vector(SS_CDEMO_SK_BUS_DATA_WIDTH-1 downto 0);
  signal cdemo_sk_inst_bus_rdat_last      : std_logic;

  signal cdemo_sk_inst_out_valid          : std_logic_vector(0 downto 0);
  signal cdemo_sk_inst_out_ready          : std_logic_vector(0 downto 0);
  signal cdemo_sk_inst_out_data           : std_logic_vector(63 downto 0);
  signal cdemo_sk_inst_out_dvalid         : std_logic_vector(0 downto 0);
  signal cdemo_sk_inst_out_last           : std_logic_vector(0 downto 0);

  signal addr_sk_inst_cmd_valid           : std_logic;
  signal addr_sk_inst_cmd_ready           : std_logic;
  signal addr_sk_inst_cmd_firstIdx        : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal addr_sk_inst_cmd_lastIdx         : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal addr_sk_inst_cmd_ctrl            : std_logic_vector(SS_ADDR_SK_BUS_ADDR_WIDTH-1 downto 0);
  signal addr_sk_inst_cmd_tag             : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal addr_sk_inst_unl_valid           : std_logic;
  signal addr_sk_inst_unl_ready           : std_logic;
  signal addr_sk_inst_unl_tag             : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal addr_sk_inst_bus_rreq_valid      : std_logic;
  signal addr_sk_inst_bus_rreq_ready      : std_logic;
  signal addr_sk_inst_bus_rreq_addr       : std_logic_vector(SS_ADDR_SK_BUS_ADDR_WIDTH-1 downto 0);
  signal addr_sk_inst_bus_rreq_len        : std_logic_vector(SS_ADDR_SK_BUS_LEN_WIDTH-1 downto 0);
  signal addr_sk_inst_bus_rdat_valid      : std_logic;
  signal addr_sk_inst_bus_rdat_ready      : std_logic;
  signal addr_sk_inst_bus_rdat_data       : std_logic_vector(SS_ADDR_SK_BUS_DATA_WIDTH-1 downto 0);
  signal addr_sk_inst_bus_rdat_last       : std_logic;

  signal addr_sk_inst_out_valid           : std_logic_vector(0 downto 0);
  signal addr_sk_inst_out_ready           : std_logic_vector(0 downto 0);
  signal addr_sk_inst_out_data            : std_logic_vector(63 downto 0);
  signal addr_sk_inst_out_dvalid          : std_logic_vector(0 downto 0);
  signal addr_sk_inst_out_last            : std_logic_vector(0 downto 0);

  signal store_sk_inst_cmd_valid          : std_logic;
  signal store_sk_inst_cmd_ready          : std_logic;
  signal store_sk_inst_cmd_firstIdx       : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal store_sk_inst_cmd_lastIdx        : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal store_sk_inst_cmd_ctrl           : std_logic_vector(SS_STORE_SK_BUS_ADDR_WIDTH-1 downto 0);
  signal store_sk_inst_cmd_tag            : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal store_sk_inst_unl_valid          : std_logic;
  signal store_sk_inst_unl_ready          : std_logic;
  signal store_sk_inst_unl_tag            : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal store_sk_inst_bus_rreq_valid     : std_logic;
  signal store_sk_inst_bus_rreq_ready     : std_logic;
  signal store_sk_inst_bus_rreq_addr      : std_logic_vector(SS_STORE_SK_BUS_ADDR_WIDTH-1 downto 0);
  signal store_sk_inst_bus_rreq_len       : std_logic_vector(SS_STORE_SK_BUS_LEN_WIDTH-1 downto 0);
  signal store_sk_inst_bus_rdat_valid     : std_logic;
  signal store_sk_inst_bus_rdat_ready     : std_logic;
  signal store_sk_inst_bus_rdat_data      : std_logic_vector(SS_STORE_SK_BUS_DATA_WIDTH-1 downto 0);
  signal store_sk_inst_bus_rdat_last      : std_logic;

  signal store_sk_inst_out_valid          : std_logic_vector(0 downto 0);
  signal store_sk_inst_out_ready          : std_logic_vector(0 downto 0);
  signal store_sk_inst_out_data           : std_logic_vector(63 downto 0);
  signal store_sk_inst_out_dvalid         : std_logic_vector(0 downto 0);
  signal store_sk_inst_out_last           : std_logic_vector(0 downto 0);

  signal quantity_inst_cmd_valid          : std_logic;
  signal quantity_inst_cmd_ready          : std_logic;
  signal quantity_inst_cmd_firstIdx       : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal quantity_inst_cmd_lastIdx        : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal quantity_inst_cmd_ctrl           : std_logic_vector(SS_QUANTITY_BUS_ADDR_WIDTH-1 downto 0);
  signal quantity_inst_cmd_tag            : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal quantity_inst_unl_valid          : std_logic;
  signal quantity_inst_unl_ready          : std_logic;
  signal quantity_inst_unl_tag            : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal quantity_inst_bus_rreq_valid     : std_logic;
  signal quantity_inst_bus_rreq_ready     : std_logic;
  signal quantity_inst_bus_rreq_addr      : std_logic_vector(SS_QUANTITY_BUS_ADDR_WIDTH-1 downto 0);
  signal quantity_inst_bus_rreq_len       : std_logic_vector(SS_QUANTITY_BUS_LEN_WIDTH-1 downto 0);
  signal quantity_inst_bus_rdat_valid     : std_logic;
  signal quantity_inst_bus_rdat_ready     : std_logic;
  signal quantity_inst_bus_rdat_data      : std_logic_vector(SS_QUANTITY_BUS_DATA_WIDTH-1 downto 0);
  signal quantity_inst_bus_rdat_last      : std_logic;

  signal quantity_inst_out_valid          : std_logic_vector(0 downto 0);
  signal quantity_inst_out_ready          : std_logic_vector(0 downto 0);
  signal quantity_inst_out_data           : std_logic_vector(63 downto 0);
  signal quantity_inst_out_dvalid         : std_logic_vector(0 downto 0);
  signal quantity_inst_out_last           : std_logic_vector(0 downto 0);

  signal sales_price_inst_cmd_valid       : std_logic;
  signal sales_price_inst_cmd_ready       : std_logic;
  signal sales_price_inst_cmd_firstIdx    : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal sales_price_inst_cmd_lastIdx     : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal sales_price_inst_cmd_ctrl        : std_logic_vector(SS_SALES_PRICE_BUS_ADDR_WIDTH-1 downto 0);
  signal sales_price_inst_cmd_tag         : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal sales_price_inst_unl_valid       : std_logic;
  signal sales_price_inst_unl_ready       : std_logic;
  signal sales_price_inst_unl_tag         : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal sales_price_inst_bus_rreq_valid  : std_logic;
  signal sales_price_inst_bus_rreq_ready  : std_logic;
  signal sales_price_inst_bus_rreq_addr   : std_logic_vector(SS_SALES_PRICE_BUS_ADDR_WIDTH-1 downto 0);
  signal sales_price_inst_bus_rreq_len    : std_logic_vector(SS_SALES_PRICE_BUS_LEN_WIDTH-1 downto 0);
  signal sales_price_inst_bus_rdat_valid  : std_logic;
  signal sales_price_inst_bus_rdat_ready  : std_logic;
  signal sales_price_inst_bus_rdat_data   : std_logic_vector(SS_SALES_PRICE_BUS_DATA_WIDTH-1 downto 0);
  signal sales_price_inst_bus_rdat_last   : std_logic;

  signal sales_price_inst_out_valid       : std_logic_vector(0 downto 0);
  signal sales_price_inst_out_ready       : std_logic_vector(0 downto 0);
  signal sales_price_inst_out_data        : std_logic_vector(63 downto 0);
  signal sales_price_inst_out_dvalid      : std_logic_vector(0 downto 0);
  signal sales_price_inst_out_last        : std_logic_vector(0 downto 0);

  signal net_profit_inst_cmd_valid        : std_logic;
  signal net_profit_inst_cmd_ready        : std_logic;
  signal net_profit_inst_cmd_firstIdx     : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal net_profit_inst_cmd_lastIdx      : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal net_profit_inst_cmd_ctrl         : std_logic_vector(SS_NET_PROFIT_BUS_ADDR_WIDTH-1 downto 0);
  signal net_profit_inst_cmd_tag          : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal net_profit_inst_unl_valid        : std_logic;
  signal net_profit_inst_unl_ready        : std_logic;
  signal net_profit_inst_unl_tag          : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal net_profit_inst_bus_rreq_valid   : std_logic;
  signal net_profit_inst_bus_rreq_ready   : std_logic;
  signal net_profit_inst_bus_rreq_addr    : std_logic_vector(SS_NET_PROFIT_BUS_ADDR_WIDTH-1 downto 0);
  signal net_profit_inst_bus_rreq_len     : std_logic_vector(SS_NET_PROFIT_BUS_LEN_WIDTH-1 downto 0);
  signal net_profit_inst_bus_rdat_valid   : std_logic;
  signal net_profit_inst_bus_rdat_ready   : std_logic;
  signal net_profit_inst_bus_rdat_data    : std_logic_vector(SS_NET_PROFIT_BUS_DATA_WIDTH-1 downto 0);
  signal net_profit_inst_bus_rdat_last    : std_logic;

  signal net_profit_inst_out_valid        : std_logic_vector(0 downto 0);
  signal net_profit_inst_out_ready        : std_logic_vector(0 downto 0);
  signal net_profit_inst_out_data         : std_logic_vector(63 downto 0);
  signal net_profit_inst_out_dvalid       : std_logic_vector(0 downto 0);
  signal net_profit_inst_out_last         : std_logic_vector(0 downto 0);

begin
  sold_date_sk_inst : ArrayReader
    generic map (
      BUS_ADDR_WIDTH     => SS_SOLD_DATE_SK_BUS_ADDR_WIDTH,
      BUS_DATA_WIDTH     => SS_SOLD_DATE_SK_BUS_DATA_WIDTH,
      BUS_LEN_WIDTH      => SS_SOLD_DATE_SK_BUS_LEN_WIDTH,
      BUS_BURST_STEP_LEN => SS_SOLD_DATE_SK_BUS_BURST_STEP_LEN,
      BUS_BURST_MAX_LEN  => SS_SOLD_DATE_SK_BUS_BURST_MAX_LEN,
      INDEX_WIDTH        => INDEX_WIDTH,
      CFG                => "prim(64)",
      CMD_TAG_ENABLE     => true,
      CMD_TAG_WIDTH      => TAG_WIDTH
    )
    port map (
      bcd_clk        => bcd_clk,
      bcd_reset      => bcd_reset,
      kcd_clk        => kcd_clk,
      kcd_reset      => kcd_reset,
      cmd_valid      => sold_date_sk_inst_cmd_valid,
      cmd_ready      => sold_date_sk_inst_cmd_ready,
      cmd_firstIdx   => sold_date_sk_inst_cmd_firstIdx,
      cmd_lastIdx    => sold_date_sk_inst_cmd_lastIdx,
      cmd_ctrl       => sold_date_sk_inst_cmd_ctrl,
      cmd_tag        => sold_date_sk_inst_cmd_tag,
      unl_valid      => sold_date_sk_inst_unl_valid,
      unl_ready      => sold_date_sk_inst_unl_ready,
      unl_tag        => sold_date_sk_inst_unl_tag,
      bus_rreq_valid => sold_date_sk_inst_bus_rreq_valid,
      bus_rreq_ready => sold_date_sk_inst_bus_rreq_ready,
      bus_rreq_addr  => sold_date_sk_inst_bus_rreq_addr,
      bus_rreq_len   => sold_date_sk_inst_bus_rreq_len,
      bus_rdat_valid => sold_date_sk_inst_bus_rdat_valid,
      bus_rdat_ready => sold_date_sk_inst_bus_rdat_ready,
      bus_rdat_data  => sold_date_sk_inst_bus_rdat_data,
      bus_rdat_last  => sold_date_sk_inst_bus_rdat_last,
      out_valid      => sold_date_sk_inst_out_valid,
      out_ready      => sold_date_sk_inst_out_ready,
      out_data       => sold_date_sk_inst_out_data,
      out_dvalid     => sold_date_sk_inst_out_dvalid,
      out_last       => sold_date_sk_inst_out_last
    );

  cdemo_sk_inst : ArrayReader
    generic map (
      BUS_ADDR_WIDTH     => SS_CDEMO_SK_BUS_ADDR_WIDTH,
      BUS_DATA_WIDTH     => SS_CDEMO_SK_BUS_DATA_WIDTH,
      BUS_LEN_WIDTH      => SS_CDEMO_SK_BUS_LEN_WIDTH,
      BUS_BURST_STEP_LEN => SS_CDEMO_SK_BUS_BURST_STEP_LEN,
      BUS_BURST_MAX_LEN  => SS_CDEMO_SK_BUS_BURST_MAX_LEN,
      INDEX_WIDTH        => INDEX_WIDTH,
      CFG                => "prim(64)",
      CMD_TAG_ENABLE     => true,
      CMD_TAG_WIDTH      => TAG_WIDTH
    )
    port map (
      bcd_clk        => bcd_clk,
      bcd_reset      => bcd_reset,
      kcd_clk        => kcd_clk,
      kcd_reset      => kcd_reset,
      cmd_valid      => cdemo_sk_inst_cmd_valid,
      cmd_ready      => cdemo_sk_inst_cmd_ready,
      cmd_firstIdx   => cdemo_sk_inst_cmd_firstIdx,
      cmd_lastIdx    => cdemo_sk_inst_cmd_lastIdx,
      cmd_ctrl       => cdemo_sk_inst_cmd_ctrl,
      cmd_tag        => cdemo_sk_inst_cmd_tag,
      unl_valid      => cdemo_sk_inst_unl_valid,
      unl_ready      => cdemo_sk_inst_unl_ready,
      unl_tag        => cdemo_sk_inst_unl_tag,
      bus_rreq_valid => cdemo_sk_inst_bus_rreq_valid,
      bus_rreq_ready => cdemo_sk_inst_bus_rreq_ready,
      bus_rreq_addr  => cdemo_sk_inst_bus_rreq_addr,
      bus_rreq_len   => cdemo_sk_inst_bus_rreq_len,
      bus_rdat_valid => cdemo_sk_inst_bus_rdat_valid,
      bus_rdat_ready => cdemo_sk_inst_bus_rdat_ready,
      bus_rdat_data  => cdemo_sk_inst_bus_rdat_data,
      bus_rdat_last  => cdemo_sk_inst_bus_rdat_last,
      out_valid      => cdemo_sk_inst_out_valid,
      out_ready      => cdemo_sk_inst_out_ready,
      out_data       => cdemo_sk_inst_out_data,
      out_dvalid     => cdemo_sk_inst_out_dvalid,
      out_last       => cdemo_sk_inst_out_last
    );

  addr_sk_inst : ArrayReader
    generic map (
      BUS_ADDR_WIDTH     => SS_ADDR_SK_BUS_ADDR_WIDTH,
      BUS_DATA_WIDTH     => SS_ADDR_SK_BUS_DATA_WIDTH,
      BUS_LEN_WIDTH      => SS_ADDR_SK_BUS_LEN_WIDTH,
      BUS_BURST_STEP_LEN => SS_ADDR_SK_BUS_BURST_STEP_LEN,
      BUS_BURST_MAX_LEN  => SS_ADDR_SK_BUS_BURST_MAX_LEN,
      INDEX_WIDTH        => INDEX_WIDTH,
      CFG                => "prim(64)",
      CMD_TAG_ENABLE     => true,
      CMD_TAG_WIDTH      => TAG_WIDTH
    )
    port map (
      bcd_clk        => bcd_clk,
      bcd_reset      => bcd_reset,
      kcd_clk        => kcd_clk,
      kcd_reset      => kcd_reset,
      cmd_valid      => addr_sk_inst_cmd_valid,
      cmd_ready      => addr_sk_inst_cmd_ready,
      cmd_firstIdx   => addr_sk_inst_cmd_firstIdx,
      cmd_lastIdx    => addr_sk_inst_cmd_lastIdx,
      cmd_ctrl       => addr_sk_inst_cmd_ctrl,
      cmd_tag        => addr_sk_inst_cmd_tag,
      unl_valid      => addr_sk_inst_unl_valid,
      unl_ready      => addr_sk_inst_unl_ready,
      unl_tag        => addr_sk_inst_unl_tag,
      bus_rreq_valid => addr_sk_inst_bus_rreq_valid,
      bus_rreq_ready => addr_sk_inst_bus_rreq_ready,
      bus_rreq_addr  => addr_sk_inst_bus_rreq_addr,
      bus_rreq_len   => addr_sk_inst_bus_rreq_len,
      bus_rdat_valid => addr_sk_inst_bus_rdat_valid,
      bus_rdat_ready => addr_sk_inst_bus_rdat_ready,
      bus_rdat_data  => addr_sk_inst_bus_rdat_data,
      bus_rdat_last  => addr_sk_inst_bus_rdat_last,
      out_valid      => addr_sk_inst_out_valid,
      out_ready      => addr_sk_inst_out_ready,
      out_data       => addr_sk_inst_out_data,
      out_dvalid     => addr_sk_inst_out_dvalid,
      out_last       => addr_sk_inst_out_last
    );

  store_sk_inst : ArrayReader
    generic map (
      BUS_ADDR_WIDTH     => SS_STORE_SK_BUS_ADDR_WIDTH,
      BUS_DATA_WIDTH     => SS_STORE_SK_BUS_DATA_WIDTH,
      BUS_LEN_WIDTH      => SS_STORE_SK_BUS_LEN_WIDTH,
      BUS_BURST_STEP_LEN => SS_STORE_SK_BUS_BURST_STEP_LEN,
      BUS_BURST_MAX_LEN  => SS_STORE_SK_BUS_BURST_MAX_LEN,
      INDEX_WIDTH        => INDEX_WIDTH,
      CFG                => "prim(64)",
      CMD_TAG_ENABLE     => true,
      CMD_TAG_WIDTH      => TAG_WIDTH
    )
    port map (
      bcd_clk        => bcd_clk,
      bcd_reset      => bcd_reset,
      kcd_clk        => kcd_clk,
      kcd_reset      => kcd_reset,
      cmd_valid      => store_sk_inst_cmd_valid,
      cmd_ready      => store_sk_inst_cmd_ready,
      cmd_firstIdx   => store_sk_inst_cmd_firstIdx,
      cmd_lastIdx    => store_sk_inst_cmd_lastIdx,
      cmd_ctrl       => store_sk_inst_cmd_ctrl,
      cmd_tag        => store_sk_inst_cmd_tag,
      unl_valid      => store_sk_inst_unl_valid,
      unl_ready      => store_sk_inst_unl_ready,
      unl_tag        => store_sk_inst_unl_tag,
      bus_rreq_valid => store_sk_inst_bus_rreq_valid,
      bus_rreq_ready => store_sk_inst_bus_rreq_ready,
      bus_rreq_addr  => store_sk_inst_bus_rreq_addr,
      bus_rreq_len   => store_sk_inst_bus_rreq_len,
      bus_rdat_valid => store_sk_inst_bus_rdat_valid,
      bus_rdat_ready => store_sk_inst_bus_rdat_ready,
      bus_rdat_data  => store_sk_inst_bus_rdat_data,
      bus_rdat_last  => store_sk_inst_bus_rdat_last,
      out_valid      => store_sk_inst_out_valid,
      out_ready      => store_sk_inst_out_ready,
      out_data       => store_sk_inst_out_data,
      out_dvalid     => store_sk_inst_out_dvalid,
      out_last       => store_sk_inst_out_last
    );

  quantity_inst : ArrayReader
    generic map (
      BUS_ADDR_WIDTH     => SS_QUANTITY_BUS_ADDR_WIDTH,
      BUS_DATA_WIDTH     => SS_QUANTITY_BUS_DATA_WIDTH,
      BUS_LEN_WIDTH      => SS_QUANTITY_BUS_LEN_WIDTH,
      BUS_BURST_STEP_LEN => SS_QUANTITY_BUS_BURST_STEP_LEN,
      BUS_BURST_MAX_LEN  => SS_QUANTITY_BUS_BURST_MAX_LEN,
      INDEX_WIDTH        => INDEX_WIDTH,
      CFG                => "prim(64)",
      CMD_TAG_ENABLE     => true,
      CMD_TAG_WIDTH      => TAG_WIDTH
    )
    port map (
      bcd_clk        => bcd_clk,
      bcd_reset      => bcd_reset,
      kcd_clk        => kcd_clk,
      kcd_reset      => kcd_reset,
      cmd_valid      => quantity_inst_cmd_valid,
      cmd_ready      => quantity_inst_cmd_ready,
      cmd_firstIdx   => quantity_inst_cmd_firstIdx,
      cmd_lastIdx    => quantity_inst_cmd_lastIdx,
      cmd_ctrl       => quantity_inst_cmd_ctrl,
      cmd_tag        => quantity_inst_cmd_tag,
      unl_valid      => quantity_inst_unl_valid,
      unl_ready      => quantity_inst_unl_ready,
      unl_tag        => quantity_inst_unl_tag,
      bus_rreq_valid => quantity_inst_bus_rreq_valid,
      bus_rreq_ready => quantity_inst_bus_rreq_ready,
      bus_rreq_addr  => quantity_inst_bus_rreq_addr,
      bus_rreq_len   => quantity_inst_bus_rreq_len,
      bus_rdat_valid => quantity_inst_bus_rdat_valid,
      bus_rdat_ready => quantity_inst_bus_rdat_ready,
      bus_rdat_data  => quantity_inst_bus_rdat_data,
      bus_rdat_last  => quantity_inst_bus_rdat_last,
      out_valid      => quantity_inst_out_valid,
      out_ready      => quantity_inst_out_ready,
      out_data       => quantity_inst_out_data,
      out_dvalid     => quantity_inst_out_dvalid,
      out_last       => quantity_inst_out_last
    );

  sales_price_inst : ArrayReader
    generic map (
      BUS_ADDR_WIDTH     => SS_SALES_PRICE_BUS_ADDR_WIDTH,
      BUS_DATA_WIDTH     => SS_SALES_PRICE_BUS_DATA_WIDTH,
      BUS_LEN_WIDTH      => SS_SALES_PRICE_BUS_LEN_WIDTH,
      BUS_BURST_STEP_LEN => SS_SALES_PRICE_BUS_BURST_STEP_LEN,
      BUS_BURST_MAX_LEN  => SS_SALES_PRICE_BUS_BURST_MAX_LEN,
      INDEX_WIDTH        => INDEX_WIDTH,
      CFG                => "prim(64)",
      CMD_TAG_ENABLE     => true,
      CMD_TAG_WIDTH      => TAG_WIDTH
    )
    port map (
      bcd_clk        => bcd_clk,
      bcd_reset      => bcd_reset,
      kcd_clk        => kcd_clk,
      kcd_reset      => kcd_reset,
      cmd_valid      => sales_price_inst_cmd_valid,
      cmd_ready      => sales_price_inst_cmd_ready,
      cmd_firstIdx   => sales_price_inst_cmd_firstIdx,
      cmd_lastIdx    => sales_price_inst_cmd_lastIdx,
      cmd_ctrl       => sales_price_inst_cmd_ctrl,
      cmd_tag        => sales_price_inst_cmd_tag,
      unl_valid      => sales_price_inst_unl_valid,
      unl_ready      => sales_price_inst_unl_ready,
      unl_tag        => sales_price_inst_unl_tag,
      bus_rreq_valid => sales_price_inst_bus_rreq_valid,
      bus_rreq_ready => sales_price_inst_bus_rreq_ready,
      bus_rreq_addr  => sales_price_inst_bus_rreq_addr,
      bus_rreq_len   => sales_price_inst_bus_rreq_len,
      bus_rdat_valid => sales_price_inst_bus_rdat_valid,
      bus_rdat_ready => sales_price_inst_bus_rdat_ready,
      bus_rdat_data  => sales_price_inst_bus_rdat_data,
      bus_rdat_last  => sales_price_inst_bus_rdat_last,
      out_valid      => sales_price_inst_out_valid,
      out_ready      => sales_price_inst_out_ready,
      out_data       => sales_price_inst_out_data,
      out_dvalid     => sales_price_inst_out_dvalid,
      out_last       => sales_price_inst_out_last
    );

  net_profit_inst : ArrayReader
    generic map (
      BUS_ADDR_WIDTH     => SS_NET_PROFIT_BUS_ADDR_WIDTH,
      BUS_DATA_WIDTH     => SS_NET_PROFIT_BUS_DATA_WIDTH,
      BUS_LEN_WIDTH      => SS_NET_PROFIT_BUS_LEN_WIDTH,
      BUS_BURST_STEP_LEN => SS_NET_PROFIT_BUS_BURST_STEP_LEN,
      BUS_BURST_MAX_LEN  => SS_NET_PROFIT_BUS_BURST_MAX_LEN,
      INDEX_WIDTH        => INDEX_WIDTH,
      CFG                => "prim(64)",
      CMD_TAG_ENABLE     => true,
      CMD_TAG_WIDTH      => TAG_WIDTH
    )
    port map (
      bcd_clk        => bcd_clk,
      bcd_reset      => bcd_reset,
      kcd_clk        => kcd_clk,
      kcd_reset      => kcd_reset,
      cmd_valid      => net_profit_inst_cmd_valid,
      cmd_ready      => net_profit_inst_cmd_ready,
      cmd_firstIdx   => net_profit_inst_cmd_firstIdx,
      cmd_lastIdx    => net_profit_inst_cmd_lastIdx,
      cmd_ctrl       => net_profit_inst_cmd_ctrl,
      cmd_tag        => net_profit_inst_cmd_tag,
      unl_valid      => net_profit_inst_unl_valid,
      unl_ready      => net_profit_inst_unl_ready,
      unl_tag        => net_profit_inst_unl_tag,
      bus_rreq_valid => net_profit_inst_bus_rreq_valid,
      bus_rreq_ready => net_profit_inst_bus_rreq_ready,
      bus_rreq_addr  => net_profit_inst_bus_rreq_addr,
      bus_rreq_len   => net_profit_inst_bus_rreq_len,
      bus_rdat_valid => net_profit_inst_bus_rdat_valid,
      bus_rdat_ready => net_profit_inst_bus_rdat_ready,
      bus_rdat_data  => net_profit_inst_bus_rdat_data,
      bus_rdat_last  => net_profit_inst_bus_rdat_last,
      out_valid      => net_profit_inst_out_valid,
      out_ready      => net_profit_inst_out_ready,
      out_data       => net_profit_inst_out_data,
      out_dvalid     => net_profit_inst_out_dvalid,
      out_last       => net_profit_inst_out_last
    );

  ss_sold_date_sk_valid            <= sold_date_sk_inst_out_valid(0);
  sold_date_sk_inst_out_ready(0)   <= ss_sold_date_sk_ready;
  ss_sold_date_sk_dvalid           <= sold_date_sk_inst_out_dvalid(0);
  ss_sold_date_sk_last             <= sold_date_sk_inst_out_last(0);
  ss_sold_date_sk                  <= sold_date_sk_inst_out_data;

  ss_sold_date_sk_bus_rreq_valid   <= sold_date_sk_inst_bus_rreq_valid;
  sold_date_sk_inst_bus_rreq_ready <= ss_sold_date_sk_bus_rreq_ready;
  ss_sold_date_sk_bus_rreq_addr    <= sold_date_sk_inst_bus_rreq_addr;
  ss_sold_date_sk_bus_rreq_len     <= sold_date_sk_inst_bus_rreq_len;
  sold_date_sk_inst_bus_rdat_valid <= ss_sold_date_sk_bus_rdat_valid;
  ss_sold_date_sk_bus_rdat_ready   <= sold_date_sk_inst_bus_rdat_ready;
  sold_date_sk_inst_bus_rdat_data  <= ss_sold_date_sk_bus_rdat_data;
  sold_date_sk_inst_bus_rdat_last  <= ss_sold_date_sk_bus_rdat_last;

  ss_sold_date_sk_unl_valid        <= sold_date_sk_inst_unl_valid;
  sold_date_sk_inst_unl_ready      <= ss_sold_date_sk_unl_ready;
  ss_sold_date_sk_unl_tag          <= sold_date_sk_inst_unl_tag;

  ss_cdemo_sk_valid                <= cdemo_sk_inst_out_valid(0);
  cdemo_sk_inst_out_ready(0)       <= ss_cdemo_sk_ready;
  ss_cdemo_sk_dvalid               <= cdemo_sk_inst_out_dvalid(0);
  ss_cdemo_sk_last                 <= cdemo_sk_inst_out_last(0);
  ss_cdemo_sk                      <= cdemo_sk_inst_out_data;

  ss_cdemo_sk_bus_rreq_valid       <= cdemo_sk_inst_bus_rreq_valid;
  cdemo_sk_inst_bus_rreq_ready     <= ss_cdemo_sk_bus_rreq_ready;
  ss_cdemo_sk_bus_rreq_addr        <= cdemo_sk_inst_bus_rreq_addr;
  ss_cdemo_sk_bus_rreq_len         <= cdemo_sk_inst_bus_rreq_len;
  cdemo_sk_inst_bus_rdat_valid     <= ss_cdemo_sk_bus_rdat_valid;
  ss_cdemo_sk_bus_rdat_ready       <= cdemo_sk_inst_bus_rdat_ready;
  cdemo_sk_inst_bus_rdat_data      <= ss_cdemo_sk_bus_rdat_data;
  cdemo_sk_inst_bus_rdat_last      <= ss_cdemo_sk_bus_rdat_last;

  ss_cdemo_sk_unl_valid            <= cdemo_sk_inst_unl_valid;
  cdemo_sk_inst_unl_ready          <= ss_cdemo_sk_unl_ready;
  ss_cdemo_sk_unl_tag              <= cdemo_sk_inst_unl_tag;

  ss_addr_sk_valid                 <= addr_sk_inst_out_valid(0);
  addr_sk_inst_out_ready(0)        <= ss_addr_sk_ready;
  ss_addr_sk_dvalid                <= addr_sk_inst_out_dvalid(0);
  ss_addr_sk_last                  <= addr_sk_inst_out_last(0);
  ss_addr_sk                       <= addr_sk_inst_out_data;

  ss_addr_sk_bus_rreq_valid        <= addr_sk_inst_bus_rreq_valid;
  addr_sk_inst_bus_rreq_ready      <= ss_addr_sk_bus_rreq_ready;
  ss_addr_sk_bus_rreq_addr         <= addr_sk_inst_bus_rreq_addr;
  ss_addr_sk_bus_rreq_len          <= addr_sk_inst_bus_rreq_len;
  addr_sk_inst_bus_rdat_valid      <= ss_addr_sk_bus_rdat_valid;
  ss_addr_sk_bus_rdat_ready        <= addr_sk_inst_bus_rdat_ready;
  addr_sk_inst_bus_rdat_data       <= ss_addr_sk_bus_rdat_data;
  addr_sk_inst_bus_rdat_last       <= ss_addr_sk_bus_rdat_last;

  ss_addr_sk_unl_valid             <= addr_sk_inst_unl_valid;
  addr_sk_inst_unl_ready           <= ss_addr_sk_unl_ready;
  ss_addr_sk_unl_tag               <= addr_sk_inst_unl_tag;

  ss_store_sk_valid                <= store_sk_inst_out_valid(0);
  store_sk_inst_out_ready(0)       <= ss_store_sk_ready;
  ss_store_sk_dvalid               <= store_sk_inst_out_dvalid(0);
  ss_store_sk_last                 <= store_sk_inst_out_last(0);
  ss_store_sk                      <= store_sk_inst_out_data;

  ss_store_sk_bus_rreq_valid       <= store_sk_inst_bus_rreq_valid;
  store_sk_inst_bus_rreq_ready     <= ss_store_sk_bus_rreq_ready;
  ss_store_sk_bus_rreq_addr        <= store_sk_inst_bus_rreq_addr;
  ss_store_sk_bus_rreq_len         <= store_sk_inst_bus_rreq_len;
  store_sk_inst_bus_rdat_valid     <= ss_store_sk_bus_rdat_valid;
  ss_store_sk_bus_rdat_ready       <= store_sk_inst_bus_rdat_ready;
  store_sk_inst_bus_rdat_data      <= ss_store_sk_bus_rdat_data;
  store_sk_inst_bus_rdat_last      <= ss_store_sk_bus_rdat_last;

  ss_store_sk_unl_valid            <= store_sk_inst_unl_valid;
  store_sk_inst_unl_ready          <= ss_store_sk_unl_ready;
  ss_store_sk_unl_tag              <= store_sk_inst_unl_tag;

  ss_quantity_valid                <= quantity_inst_out_valid(0);
  quantity_inst_out_ready(0)       <= ss_quantity_ready;
  ss_quantity_dvalid               <= quantity_inst_out_dvalid(0);
  ss_quantity_last                 <= quantity_inst_out_last(0);
  ss_quantity                      <= quantity_inst_out_data;

  ss_quantity_bus_rreq_valid       <= quantity_inst_bus_rreq_valid;
  quantity_inst_bus_rreq_ready     <= ss_quantity_bus_rreq_ready;
  ss_quantity_bus_rreq_addr        <= quantity_inst_bus_rreq_addr;
  ss_quantity_bus_rreq_len         <= quantity_inst_bus_rreq_len;
  quantity_inst_bus_rdat_valid     <= ss_quantity_bus_rdat_valid;
  ss_quantity_bus_rdat_ready       <= quantity_inst_bus_rdat_ready;
  quantity_inst_bus_rdat_data      <= ss_quantity_bus_rdat_data;
  quantity_inst_bus_rdat_last      <= ss_quantity_bus_rdat_last;

  ss_quantity_unl_valid            <= quantity_inst_unl_valid;
  quantity_inst_unl_ready          <= ss_quantity_unl_ready;
  ss_quantity_unl_tag              <= quantity_inst_unl_tag;

  ss_sales_price_valid             <= sales_price_inst_out_valid(0);
  sales_price_inst_out_ready(0)    <= ss_sales_price_ready;
  ss_sales_price_dvalid            <= sales_price_inst_out_dvalid(0);
  ss_sales_price_last              <= sales_price_inst_out_last(0);
  ss_sales_price                   <= sales_price_inst_out_data;

  ss_sales_price_bus_rreq_valid    <= sales_price_inst_bus_rreq_valid;
  sales_price_inst_bus_rreq_ready  <= ss_sales_price_bus_rreq_ready;
  ss_sales_price_bus_rreq_addr     <= sales_price_inst_bus_rreq_addr;
  ss_sales_price_bus_rreq_len      <= sales_price_inst_bus_rreq_len;
  sales_price_inst_bus_rdat_valid  <= ss_sales_price_bus_rdat_valid;
  ss_sales_price_bus_rdat_ready    <= sales_price_inst_bus_rdat_ready;
  sales_price_inst_bus_rdat_data   <= ss_sales_price_bus_rdat_data;
  sales_price_inst_bus_rdat_last   <= ss_sales_price_bus_rdat_last;

  ss_sales_price_unl_valid         <= sales_price_inst_unl_valid;
  sales_price_inst_unl_ready       <= ss_sales_price_unl_ready;
  ss_sales_price_unl_tag           <= sales_price_inst_unl_tag;

  ss_net_profit_valid              <= net_profit_inst_out_valid(0);
  net_profit_inst_out_ready(0)     <= ss_net_profit_ready;
  ss_net_profit_dvalid             <= net_profit_inst_out_dvalid(0);
  ss_net_profit_last               <= net_profit_inst_out_last(0);
  ss_net_profit                    <= net_profit_inst_out_data;

  ss_net_profit_bus_rreq_valid     <= net_profit_inst_bus_rreq_valid;
  net_profit_inst_bus_rreq_ready   <= ss_net_profit_bus_rreq_ready;
  ss_net_profit_bus_rreq_addr      <= net_profit_inst_bus_rreq_addr;
  ss_net_profit_bus_rreq_len       <= net_profit_inst_bus_rreq_len;
  net_profit_inst_bus_rdat_valid   <= ss_net_profit_bus_rdat_valid;
  ss_net_profit_bus_rdat_ready     <= net_profit_inst_bus_rdat_ready;
  net_profit_inst_bus_rdat_data    <= ss_net_profit_bus_rdat_data;
  net_profit_inst_bus_rdat_last    <= ss_net_profit_bus_rdat_last;

  ss_net_profit_unl_valid          <= net_profit_inst_unl_valid;
  net_profit_inst_unl_ready        <= ss_net_profit_unl_ready;
  ss_net_profit_unl_tag            <= net_profit_inst_unl_tag;

  sold_date_sk_inst_cmd_valid    <= ss_sold_date_sk_cmd_valid;
  ss_sold_date_sk_cmd_ready      <= sold_date_sk_inst_cmd_ready;
  sold_date_sk_inst_cmd_firstIdx <= ss_sold_date_sk_cmd_firstIdx;
  sold_date_sk_inst_cmd_lastIdx  <= ss_sold_date_sk_cmd_lastIdx;
  sold_date_sk_inst_cmd_ctrl     <= ss_sold_date_sk_cmd_ctrl;
  sold_date_sk_inst_cmd_tag      <= ss_sold_date_sk_cmd_tag;

  cdemo_sk_inst_cmd_valid        <= ss_cdemo_sk_cmd_valid;
  ss_cdemo_sk_cmd_ready          <= cdemo_sk_inst_cmd_ready;
  cdemo_sk_inst_cmd_firstIdx     <= ss_cdemo_sk_cmd_firstIdx;
  cdemo_sk_inst_cmd_lastIdx      <= ss_cdemo_sk_cmd_lastIdx;
  cdemo_sk_inst_cmd_ctrl         <= ss_cdemo_sk_cmd_ctrl;
  cdemo_sk_inst_cmd_tag          <= ss_cdemo_sk_cmd_tag;

  addr_sk_inst_cmd_valid         <= ss_addr_sk_cmd_valid;
  ss_addr_sk_cmd_ready           <= addr_sk_inst_cmd_ready;
  addr_sk_inst_cmd_firstIdx      <= ss_addr_sk_cmd_firstIdx;
  addr_sk_inst_cmd_lastIdx       <= ss_addr_sk_cmd_lastIdx;
  addr_sk_inst_cmd_ctrl          <= ss_addr_sk_cmd_ctrl;
  addr_sk_inst_cmd_tag           <= ss_addr_sk_cmd_tag;

  store_sk_inst_cmd_valid        <= ss_store_sk_cmd_valid;
  ss_store_sk_cmd_ready          <= store_sk_inst_cmd_ready;
  store_sk_inst_cmd_firstIdx     <= ss_store_sk_cmd_firstIdx;
  store_sk_inst_cmd_lastIdx      <= ss_store_sk_cmd_lastIdx;
  store_sk_inst_cmd_ctrl         <= ss_store_sk_cmd_ctrl;
  store_sk_inst_cmd_tag          <= ss_store_sk_cmd_tag;

  quantity_inst_cmd_valid        <= ss_quantity_cmd_valid;
  ss_quantity_cmd_ready          <= quantity_inst_cmd_ready;
  quantity_inst_cmd_firstIdx     <= ss_quantity_cmd_firstIdx;
  quantity_inst_cmd_lastIdx      <= ss_quantity_cmd_lastIdx;
  quantity_inst_cmd_ctrl         <= ss_quantity_cmd_ctrl;
  quantity_inst_cmd_tag          <= ss_quantity_cmd_tag;

  sales_price_inst_cmd_valid     <= ss_sales_price_cmd_valid;
  ss_sales_price_cmd_ready       <= sales_price_inst_cmd_ready;
  sales_price_inst_cmd_firstIdx  <= ss_sales_price_cmd_firstIdx;
  sales_price_inst_cmd_lastIdx   <= ss_sales_price_cmd_lastIdx;
  sales_price_inst_cmd_ctrl      <= ss_sales_price_cmd_ctrl;
  sales_price_inst_cmd_tag       <= ss_sales_price_cmd_tag;

  net_profit_inst_cmd_valid      <= ss_net_profit_cmd_valid;
  ss_net_profit_cmd_ready        <= net_profit_inst_cmd_ready;
  net_profit_inst_cmd_firstIdx   <= ss_net_profit_cmd_firstIdx;
  net_profit_inst_cmd_lastIdx    <= ss_net_profit_cmd_lastIdx;
  net_profit_inst_cmd_ctrl       <= ss_net_profit_cmd_ctrl;
  net_profit_inst_cmd_tag        <= ss_net_profit_cmd_tag;

end architecture;
