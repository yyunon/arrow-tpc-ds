-- Copyright 2018-2019 Delft University of Technology
--
-- Licensed under the Apache License, Version 2.0 (the "License");
-- you may not use this file except in compliance with the License.
-- You may obtain a copy of the License at
--
--     http://www.apache.org/licenses/LICENSE-2.0
--
-- Unless required by applicable law or agreed to in writing, software
-- distributed under the License is distributed on an "AS IS" BASIS,
-- WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
-- See the License for the specific language governing permissions and
-- limitations under the License.
--
-- This file was generated by Fletchgen. Modify this file at your own risk.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library work;
use work.Array_pkg.all;
use work.mmio_pkg.all;

entity Join_Nucleus is
  generic (
    INDEX_WIDTH                    : integer := 32;
    TAG_WIDTH                      : integer := 1;
    SS_SOLD_DATE_SK_BUS_ADDR_WIDTH : integer := 64;
    SS_CDEMO_SK_BUS_ADDR_WIDTH     : integer := 64;
    SS_ADDR_SK_BUS_ADDR_WIDTH      : integer := 64;
    SS_STORE_SK_BUS_ADDR_WIDTH     : integer := 64;
    SS_QUANTITY_BUS_ADDR_WIDTH     : integer := 64;
    SS_SALES_PRICE_BUS_ADDR_WIDTH  : integer := 64;
    SS_NET_PROFIT_BUS_ADDR_WIDTH   : integer := 64
  );
  port (
    kcd_clk                      : in  std_logic;
    kcd_reset                    : in  std_logic;
    mmio_awvalid                 : in  std_logic;
    mmio_awready                 : out std_logic;
    mmio_awaddr                  : in  std_logic_vector(31 downto 0);
    mmio_wvalid                  : in  std_logic;
    mmio_wready                  : out std_logic;
    mmio_wdata                   : in  std_logic_vector(31 downto 0);
    mmio_wstrb                   : in  std_logic_vector(3 downto 0);
    mmio_bvalid                  : out std_logic;
    mmio_bready                  : in  std_logic;
    mmio_bresp                   : out std_logic_vector(1 downto 0);
    mmio_arvalid                 : in  std_logic;
    mmio_arready                 : out std_logic;
    mmio_araddr                  : in  std_logic_vector(31 downto 0);
    mmio_rvalid                  : out std_logic;
    mmio_rready                  : in  std_logic;
    mmio_rdata                   : out std_logic_vector(31 downto 0);
    mmio_rresp                   : out std_logic_vector(1 downto 0);
    ss_sold_date_sk_valid        : in  std_logic;
    ss_sold_date_sk_ready        : out std_logic;
    ss_sold_date_sk_dvalid       : in  std_logic;
    ss_sold_date_sk_last         : in  std_logic;
    ss_sold_date_sk              : in  std_logic_vector(63 downto 0);
    ss_cdemo_sk_valid            : in  std_logic;
    ss_cdemo_sk_ready            : out std_logic;
    ss_cdemo_sk_dvalid           : in  std_logic;
    ss_cdemo_sk_last             : in  std_logic;
    ss_cdemo_sk                  : in  std_logic_vector(63 downto 0);
    ss_addr_sk_valid             : in  std_logic;
    ss_addr_sk_ready             : out std_logic;
    ss_addr_sk_dvalid            : in  std_logic;
    ss_addr_sk_last              : in  std_logic;
    ss_addr_sk                   : in  std_logic_vector(63 downto 0);
    ss_store_sk_valid            : in  std_logic;
    ss_store_sk_ready            : out std_logic;
    ss_store_sk_dvalid           : in  std_logic;
    ss_store_sk_last             : in  std_logic;
    ss_store_sk                  : in  std_logic_vector(63 downto 0);
    ss_quantity_valid            : in  std_logic;
    ss_quantity_ready            : out std_logic;
    ss_quantity_dvalid           : in  std_logic;
    ss_quantity_last             : in  std_logic;
    ss_quantity                  : in  std_logic_vector(63 downto 0);
    ss_sales_price_valid         : in  std_logic;
    ss_sales_price_ready         : out std_logic;
    ss_sales_price_dvalid        : in  std_logic;
    ss_sales_price_last          : in  std_logic;
    ss_sales_price               : in  std_logic_vector(63 downto 0);
    ss_net_profit_valid          : in  std_logic;
    ss_net_profit_ready          : out std_logic;
    ss_net_profit_dvalid         : in  std_logic;
    ss_net_profit_last           : in  std_logic;
    ss_net_profit                : in  std_logic_vector(63 downto 0);
    ss_sold_date_sk_unl_valid    : in  std_logic;
    ss_sold_date_sk_unl_ready    : out std_logic;
    ss_sold_date_sk_unl_tag      : in  std_logic_vector(TAG_WIDTH-1 downto 0);
    ss_cdemo_sk_unl_valid        : in  std_logic;
    ss_cdemo_sk_unl_ready        : out std_logic;
    ss_cdemo_sk_unl_tag          : in  std_logic_vector(TAG_WIDTH-1 downto 0);
    ss_addr_sk_unl_valid         : in  std_logic;
    ss_addr_sk_unl_ready         : out std_logic;
    ss_addr_sk_unl_tag           : in  std_logic_vector(TAG_WIDTH-1 downto 0);
    ss_store_sk_unl_valid        : in  std_logic;
    ss_store_sk_unl_ready        : out std_logic;
    ss_store_sk_unl_tag          : in  std_logic_vector(TAG_WIDTH-1 downto 0);
    ss_quantity_unl_valid        : in  std_logic;
    ss_quantity_unl_ready        : out std_logic;
    ss_quantity_unl_tag          : in  std_logic_vector(TAG_WIDTH-1 downto 0);
    ss_sales_price_unl_valid     : in  std_logic;
    ss_sales_price_unl_ready     : out std_logic;
    ss_sales_price_unl_tag       : in  std_logic_vector(TAG_WIDTH-1 downto 0);
    ss_net_profit_unl_valid      : in  std_logic;
    ss_net_profit_unl_ready      : out std_logic;
    ss_net_profit_unl_tag        : in  std_logic_vector(TAG_WIDTH-1 downto 0);
    ss_sold_date_sk_cmd_valid    : out std_logic;
    ss_sold_date_sk_cmd_ready    : in  std_logic;
    ss_sold_date_sk_cmd_firstIdx : out std_logic_vector(INDEX_WIDTH-1 downto 0);
    ss_sold_date_sk_cmd_lastIdx  : out std_logic_vector(INDEX_WIDTH-1 downto 0);
    ss_sold_date_sk_cmd_ctrl     : out std_logic_vector(SS_SOLD_DATE_SK_BUS_ADDR_WIDTH-1 downto 0);
    ss_sold_date_sk_cmd_tag      : out std_logic_vector(TAG_WIDTH-1 downto 0);
    ss_cdemo_sk_cmd_valid        : out std_logic;
    ss_cdemo_sk_cmd_ready        : in  std_logic;
    ss_cdemo_sk_cmd_firstIdx     : out std_logic_vector(INDEX_WIDTH-1 downto 0);
    ss_cdemo_sk_cmd_lastIdx      : out std_logic_vector(INDEX_WIDTH-1 downto 0);
    ss_cdemo_sk_cmd_ctrl         : out std_logic_vector(SS_CDEMO_SK_BUS_ADDR_WIDTH-1 downto 0);
    ss_cdemo_sk_cmd_tag          : out std_logic_vector(TAG_WIDTH-1 downto 0);
    ss_addr_sk_cmd_valid         : out std_logic;
    ss_addr_sk_cmd_ready         : in  std_logic;
    ss_addr_sk_cmd_firstIdx      : out std_logic_vector(INDEX_WIDTH-1 downto 0);
    ss_addr_sk_cmd_lastIdx       : out std_logic_vector(INDEX_WIDTH-1 downto 0);
    ss_addr_sk_cmd_ctrl          : out std_logic_vector(SS_ADDR_SK_BUS_ADDR_WIDTH-1 downto 0);
    ss_addr_sk_cmd_tag           : out std_logic_vector(TAG_WIDTH-1 downto 0);
    ss_store_sk_cmd_valid        : out std_logic;
    ss_store_sk_cmd_ready        : in  std_logic;
    ss_store_sk_cmd_firstIdx     : out std_logic_vector(INDEX_WIDTH-1 downto 0);
    ss_store_sk_cmd_lastIdx      : out std_logic_vector(INDEX_WIDTH-1 downto 0);
    ss_store_sk_cmd_ctrl         : out std_logic_vector(SS_STORE_SK_BUS_ADDR_WIDTH-1 downto 0);
    ss_store_sk_cmd_tag          : out std_logic_vector(TAG_WIDTH-1 downto 0);
    ss_quantity_cmd_valid        : out std_logic;
    ss_quantity_cmd_ready        : in  std_logic;
    ss_quantity_cmd_firstIdx     : out std_logic_vector(INDEX_WIDTH-1 downto 0);
    ss_quantity_cmd_lastIdx      : out std_logic_vector(INDEX_WIDTH-1 downto 0);
    ss_quantity_cmd_ctrl         : out std_logic_vector(SS_QUANTITY_BUS_ADDR_WIDTH-1 downto 0);
    ss_quantity_cmd_tag          : out std_logic_vector(TAG_WIDTH-1 downto 0);
    ss_sales_price_cmd_valid     : out std_logic;
    ss_sales_price_cmd_ready     : in  std_logic;
    ss_sales_price_cmd_firstIdx  : out std_logic_vector(INDEX_WIDTH-1 downto 0);
    ss_sales_price_cmd_lastIdx   : out std_logic_vector(INDEX_WIDTH-1 downto 0);
    ss_sales_price_cmd_ctrl      : out std_logic_vector(SS_SALES_PRICE_BUS_ADDR_WIDTH-1 downto 0);
    ss_sales_price_cmd_tag       : out std_logic_vector(TAG_WIDTH-1 downto 0);
    ss_net_profit_cmd_valid      : out std_logic;
    ss_net_profit_cmd_ready      : in  std_logic;
    ss_net_profit_cmd_firstIdx   : out std_logic_vector(INDEX_WIDTH-1 downto 0);
    ss_net_profit_cmd_lastIdx    : out std_logic_vector(INDEX_WIDTH-1 downto 0);
    ss_net_profit_cmd_ctrl       : out std_logic_vector(SS_NET_PROFIT_BUS_ADDR_WIDTH-1 downto 0);
    ss_net_profit_cmd_tag        : out std_logic_vector(TAG_WIDTH-1 downto 0)
  );
end entity;

architecture Implementation of Join_Nucleus is
  component Join is
    generic (
      INDEX_WIDTH : integer := 32;
      TAG_WIDTH   : integer := 1
    );
    port (
      kcd_clk                      : in  std_logic;
      kcd_reset                    : in  std_logic;
      ss_sold_date_sk_valid        : in  std_logic;
      ss_sold_date_sk_ready        : out std_logic;
      ss_sold_date_sk_dvalid       : in  std_logic;
      ss_sold_date_sk_last         : in  std_logic;
      ss_sold_date_sk              : in  std_logic_vector(63 downto 0);
      ss_cdemo_sk_valid            : in  std_logic;
      ss_cdemo_sk_ready            : out std_logic;
      ss_cdemo_sk_dvalid           : in  std_logic;
      ss_cdemo_sk_last             : in  std_logic;
      ss_cdemo_sk                  : in  std_logic_vector(63 downto 0);
      ss_addr_sk_valid             : in  std_logic;
      ss_addr_sk_ready             : out std_logic;
      ss_addr_sk_dvalid            : in  std_logic;
      ss_addr_sk_last              : in  std_logic;
      ss_addr_sk                   : in  std_logic_vector(63 downto 0);
      ss_store_sk_valid            : in  std_logic;
      ss_store_sk_ready            : out std_logic;
      ss_store_sk_dvalid           : in  std_logic;
      ss_store_sk_last             : in  std_logic;
      ss_store_sk                  : in  std_logic_vector(63 downto 0);
      ss_quantity_valid            : in  std_logic;
      ss_quantity_ready            : out std_logic;
      ss_quantity_dvalid           : in  std_logic;
      ss_quantity_last             : in  std_logic;
      ss_quantity                  : in  std_logic_vector(63 downto 0);
      ss_sales_price_valid         : in  std_logic;
      ss_sales_price_ready         : out std_logic;
      ss_sales_price_dvalid        : in  std_logic;
      ss_sales_price_last          : in  std_logic;
      ss_sales_price               : in  std_logic_vector(63 downto 0);
      ss_net_profit_valid          : in  std_logic;
      ss_net_profit_ready          : out std_logic;
      ss_net_profit_dvalid         : in  std_logic;
      ss_net_profit_last           : in  std_logic;
      ss_net_profit                : in  std_logic_vector(63 downto 0);
      ss_sold_date_sk_unl_valid    : in  std_logic;
      ss_sold_date_sk_unl_ready    : out std_logic;
      ss_sold_date_sk_unl_tag      : in  std_logic_vector(TAG_WIDTH-1 downto 0);
      ss_cdemo_sk_unl_valid        : in  std_logic;
      ss_cdemo_sk_unl_ready        : out std_logic;
      ss_cdemo_sk_unl_tag          : in  std_logic_vector(TAG_WIDTH-1 downto 0);
      ss_addr_sk_unl_valid         : in  std_logic;
      ss_addr_sk_unl_ready         : out std_logic;
      ss_addr_sk_unl_tag           : in  std_logic_vector(TAG_WIDTH-1 downto 0);
      ss_store_sk_unl_valid        : in  std_logic;
      ss_store_sk_unl_ready        : out std_logic;
      ss_store_sk_unl_tag          : in  std_logic_vector(TAG_WIDTH-1 downto 0);
      ss_quantity_unl_valid        : in  std_logic;
      ss_quantity_unl_ready        : out std_logic;
      ss_quantity_unl_tag          : in  std_logic_vector(TAG_WIDTH-1 downto 0);
      ss_sales_price_unl_valid     : in  std_logic;
      ss_sales_price_unl_ready     : out std_logic;
      ss_sales_price_unl_tag       : in  std_logic_vector(TAG_WIDTH-1 downto 0);
      ss_net_profit_unl_valid      : in  std_logic;
      ss_net_profit_unl_ready      : out std_logic;
      ss_net_profit_unl_tag        : in  std_logic_vector(TAG_WIDTH-1 downto 0);
      ss_sold_date_sk_cmd_valid    : out std_logic;
      ss_sold_date_sk_cmd_ready    : in  std_logic;
      ss_sold_date_sk_cmd_firstIdx : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      ss_sold_date_sk_cmd_lastIdx  : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      ss_sold_date_sk_cmd_tag      : out std_logic_vector(TAG_WIDTH-1 downto 0);
      ss_cdemo_sk_cmd_valid        : out std_logic;
      ss_cdemo_sk_cmd_ready        : in  std_logic;
      ss_cdemo_sk_cmd_firstIdx     : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      ss_cdemo_sk_cmd_lastIdx      : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      ss_cdemo_sk_cmd_tag          : out std_logic_vector(TAG_WIDTH-1 downto 0);
      ss_addr_sk_cmd_valid         : out std_logic;
      ss_addr_sk_cmd_ready         : in  std_logic;
      ss_addr_sk_cmd_firstIdx      : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      ss_addr_sk_cmd_lastIdx       : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      ss_addr_sk_cmd_tag           : out std_logic_vector(TAG_WIDTH-1 downto 0);
      ss_store_sk_cmd_valid        : out std_logic;
      ss_store_sk_cmd_ready        : in  std_logic;
      ss_store_sk_cmd_firstIdx     : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      ss_store_sk_cmd_lastIdx      : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      ss_store_sk_cmd_tag          : out std_logic_vector(TAG_WIDTH-1 downto 0);
      ss_quantity_cmd_valid        : out std_logic;
      ss_quantity_cmd_ready        : in  std_logic;
      ss_quantity_cmd_firstIdx     : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      ss_quantity_cmd_lastIdx      : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      ss_quantity_cmd_tag          : out std_logic_vector(TAG_WIDTH-1 downto 0);
      ss_sales_price_cmd_valid     : out std_logic;
      ss_sales_price_cmd_ready     : in  std_logic;
      ss_sales_price_cmd_firstIdx  : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      ss_sales_price_cmd_lastIdx   : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      ss_sales_price_cmd_tag       : out std_logic_vector(TAG_WIDTH-1 downto 0);
      ss_net_profit_cmd_valid      : out std_logic;
      ss_net_profit_cmd_ready      : in  std_logic;
      ss_net_profit_cmd_firstIdx   : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      ss_net_profit_cmd_lastIdx    : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      ss_net_profit_cmd_tag        : out std_logic_vector(TAG_WIDTH-1 downto 0);
      start                        : in  std_logic;
      stop                         : in  std_logic;
      reset                        : in  std_logic;
      idle                         : out std_logic;
      busy                         : out std_logic;
      done                         : out std_logic;
      result                       : out std_logic_vector(63 downto 0);
      ss_firstidx                  : in  std_logic_vector(31 downto 0);
      ss_lastidx                   : in  std_logic_vector(31 downto 0)
    );
  end component;

  signal Join_inst_ss_sold_date_sk_valid                    : std_logic;
  signal Join_inst_ss_sold_date_sk_ready                    : std_logic;
  signal Join_inst_ss_sold_date_sk_dvalid                   : std_logic;
  signal Join_inst_ss_sold_date_sk_last                     : std_logic;
  signal Join_inst_ss_sold_date_sk                          : std_logic_vector(63 downto 0);

  signal Join_inst_ss_cdemo_sk_valid                        : std_logic;
  signal Join_inst_ss_cdemo_sk_ready                        : std_logic;
  signal Join_inst_ss_cdemo_sk_dvalid                       : std_logic;
  signal Join_inst_ss_cdemo_sk_last                         : std_logic;
  signal Join_inst_ss_cdemo_sk                              : std_logic_vector(63 downto 0);

  signal Join_inst_ss_addr_sk_valid                         : std_logic;
  signal Join_inst_ss_addr_sk_ready                         : std_logic;
  signal Join_inst_ss_addr_sk_dvalid                        : std_logic;
  signal Join_inst_ss_addr_sk_last                          : std_logic;
  signal Join_inst_ss_addr_sk                               : std_logic_vector(63 downto 0);

  signal Join_inst_ss_store_sk_valid                        : std_logic;
  signal Join_inst_ss_store_sk_ready                        : std_logic;
  signal Join_inst_ss_store_sk_dvalid                       : std_logic;
  signal Join_inst_ss_store_sk_last                         : std_logic;
  signal Join_inst_ss_store_sk                              : std_logic_vector(63 downto 0);

  signal Join_inst_ss_quantity_valid                        : std_logic;
  signal Join_inst_ss_quantity_ready                        : std_logic;
  signal Join_inst_ss_quantity_dvalid                       : std_logic;
  signal Join_inst_ss_quantity_last                         : std_logic;
  signal Join_inst_ss_quantity                              : std_logic_vector(63 downto 0);

  signal Join_inst_ss_sales_price_valid                     : std_logic;
  signal Join_inst_ss_sales_price_ready                     : std_logic;
  signal Join_inst_ss_sales_price_dvalid                    : std_logic;
  signal Join_inst_ss_sales_price_last                      : std_logic;
  signal Join_inst_ss_sales_price                           : std_logic_vector(63 downto 0);

  signal Join_inst_ss_net_profit_valid                      : std_logic;
  signal Join_inst_ss_net_profit_ready                      : std_logic;
  signal Join_inst_ss_net_profit_dvalid                     : std_logic;
  signal Join_inst_ss_net_profit_last                       : std_logic;
  signal Join_inst_ss_net_profit                            : std_logic_vector(63 downto 0);

  signal Join_inst_ss_sold_date_sk_unl_valid                : std_logic;
  signal Join_inst_ss_sold_date_sk_unl_ready                : std_logic;
  signal Join_inst_ss_sold_date_sk_unl_tag                  : std_logic_vector(0 downto 0);

  signal Join_inst_ss_cdemo_sk_unl_valid                    : std_logic;
  signal Join_inst_ss_cdemo_sk_unl_ready                    : std_logic;
  signal Join_inst_ss_cdemo_sk_unl_tag                      : std_logic_vector(0 downto 0);

  signal Join_inst_ss_addr_sk_unl_valid                     : std_logic;
  signal Join_inst_ss_addr_sk_unl_ready                     : std_logic;
  signal Join_inst_ss_addr_sk_unl_tag                       : std_logic_vector(0 downto 0);

  signal Join_inst_ss_store_sk_unl_valid                    : std_logic;
  signal Join_inst_ss_store_sk_unl_ready                    : std_logic;
  signal Join_inst_ss_store_sk_unl_tag                      : std_logic_vector(0 downto 0);

  signal Join_inst_ss_quantity_unl_valid                    : std_logic;
  signal Join_inst_ss_quantity_unl_ready                    : std_logic;
  signal Join_inst_ss_quantity_unl_tag                      : std_logic_vector(0 downto 0);

  signal Join_inst_ss_sales_price_unl_valid                 : std_logic;
  signal Join_inst_ss_sales_price_unl_ready                 : std_logic;
  signal Join_inst_ss_sales_price_unl_tag                   : std_logic_vector(0 downto 0);

  signal Join_inst_ss_net_profit_unl_valid                  : std_logic;
  signal Join_inst_ss_net_profit_unl_ready                  : std_logic;
  signal Join_inst_ss_net_profit_unl_tag                    : std_logic_vector(0 downto 0);

  signal Join_inst_ss_sold_date_sk_cmd_valid                : std_logic;
  signal Join_inst_ss_sold_date_sk_cmd_ready                : std_logic;
  signal Join_inst_ss_sold_date_sk_cmd_firstIdx             : std_logic_vector(31 downto 0);
  signal Join_inst_ss_sold_date_sk_cmd_lastIdx              : std_logic_vector(31 downto 0);
  signal Join_inst_ss_sold_date_sk_cmd_tag                  : std_logic_vector(0 downto 0);

  signal Join_inst_ss_cdemo_sk_cmd_valid                    : std_logic;
  signal Join_inst_ss_cdemo_sk_cmd_ready                    : std_logic;
  signal Join_inst_ss_cdemo_sk_cmd_firstIdx                 : std_logic_vector(31 downto 0);
  signal Join_inst_ss_cdemo_sk_cmd_lastIdx                  : std_logic_vector(31 downto 0);
  signal Join_inst_ss_cdemo_sk_cmd_tag                      : std_logic_vector(0 downto 0);

  signal Join_inst_ss_addr_sk_cmd_valid                     : std_logic;
  signal Join_inst_ss_addr_sk_cmd_ready                     : std_logic;
  signal Join_inst_ss_addr_sk_cmd_firstIdx                  : std_logic_vector(31 downto 0);
  signal Join_inst_ss_addr_sk_cmd_lastIdx                   : std_logic_vector(31 downto 0);
  signal Join_inst_ss_addr_sk_cmd_tag                       : std_logic_vector(0 downto 0);

  signal Join_inst_ss_store_sk_cmd_valid                    : std_logic;
  signal Join_inst_ss_store_sk_cmd_ready                    : std_logic;
  signal Join_inst_ss_store_sk_cmd_firstIdx                 : std_logic_vector(31 downto 0);
  signal Join_inst_ss_store_sk_cmd_lastIdx                  : std_logic_vector(31 downto 0);
  signal Join_inst_ss_store_sk_cmd_tag                      : std_logic_vector(0 downto 0);

  signal Join_inst_ss_quantity_cmd_valid                    : std_logic;
  signal Join_inst_ss_quantity_cmd_ready                    : std_logic;
  signal Join_inst_ss_quantity_cmd_firstIdx                 : std_logic_vector(31 downto 0);
  signal Join_inst_ss_quantity_cmd_lastIdx                  : std_logic_vector(31 downto 0);
  signal Join_inst_ss_quantity_cmd_tag                      : std_logic_vector(0 downto 0);

  signal Join_inst_ss_sales_price_cmd_valid                 : std_logic;
  signal Join_inst_ss_sales_price_cmd_ready                 : std_logic;
  signal Join_inst_ss_sales_price_cmd_firstIdx              : std_logic_vector(31 downto 0);
  signal Join_inst_ss_sales_price_cmd_lastIdx               : std_logic_vector(31 downto 0);
  signal Join_inst_ss_sales_price_cmd_tag                   : std_logic_vector(0 downto 0);

  signal Join_inst_ss_net_profit_cmd_valid                  : std_logic;
  signal Join_inst_ss_net_profit_cmd_ready                  : std_logic;
  signal Join_inst_ss_net_profit_cmd_firstIdx               : std_logic_vector(31 downto 0);
  signal Join_inst_ss_net_profit_cmd_lastIdx                : std_logic_vector(31 downto 0);
  signal Join_inst_ss_net_profit_cmd_tag                    : std_logic_vector(0 downto 0);

  signal Join_inst_start                                    : std_logic;
  signal Join_inst_stop                                     : std_logic;
  signal Join_inst_reset                                    : std_logic;
  signal Join_inst_idle                                     : std_logic;
  signal Join_inst_busy                                     : std_logic;
  signal Join_inst_done                                     : std_logic;
  signal Join_inst_result                                   : std_logic_vector(63 downto 0);
  signal Join_inst_ss_firstidx                              : std_logic_vector(31 downto 0);
  signal Join_inst_ss_lastidx                               : std_logic_vector(31 downto 0);
  signal mmio_inst_f_start_data                             : std_logic;
  signal mmio_inst_f_stop_data                              : std_logic;
  signal mmio_inst_f_reset_data                             : std_logic;
  signal mmio_inst_f_idle_write_data                        : std_logic;
  signal mmio_inst_f_busy_write_data                        : std_logic;
  signal mmio_inst_f_done_write_data                        : std_logic;
  signal mmio_inst_f_result_write_data                      : std_logic_vector(63 downto 0);
  signal mmio_inst_f_ss_firstidx_data                       : std_logic_vector(31 downto 0);
  signal mmio_inst_f_ss_lastidx_data                        : std_logic_vector(31 downto 0);
  signal mmio_inst_f_ss_sold_date_sk_values_data            : std_logic_vector(63 downto 0);
  signal mmio_inst_f_ss_cdemo_sk_values_data                : std_logic_vector(63 downto 0);
  signal mmio_inst_f_ss_addr_sk_values_data                 : std_logic_vector(63 downto 0);
  signal mmio_inst_f_ss_store_sk_values_data                : std_logic_vector(63 downto 0);
  signal mmio_inst_f_ss_quantity_values_data                : std_logic_vector(63 downto 0);
  signal mmio_inst_f_ss_sales_price_values_data             : std_logic_vector(63 downto 0);
  signal mmio_inst_f_ss_net_profit_values_data              : std_logic_vector(63 downto 0);
  signal mmio_inst_f_Profile_enable_data                    : std_logic;
  signal mmio_inst_f_Profile_clear_data                     : std_logic;
  signal mmio_inst_mmio_awvalid                             : std_logic;
  signal mmio_inst_mmio_awready                             : std_logic;
  signal mmio_inst_mmio_awaddr                              : std_logic_vector(31 downto 0);
  signal mmio_inst_mmio_wvalid                              : std_logic;
  signal mmio_inst_mmio_wready                              : std_logic;
  signal mmio_inst_mmio_wdata                               : std_logic_vector(31 downto 0);
  signal mmio_inst_mmio_wstrb                               : std_logic_vector(3 downto 0);
  signal mmio_inst_mmio_bvalid                              : std_logic;
  signal mmio_inst_mmio_bready                              : std_logic;
  signal mmio_inst_mmio_bresp                               : std_logic_vector(1 downto 0);
  signal mmio_inst_mmio_arvalid                             : std_logic;
  signal mmio_inst_mmio_arready                             : std_logic;
  signal mmio_inst_mmio_araddr                              : std_logic_vector(31 downto 0);
  signal mmio_inst_mmio_rvalid                              : std_logic;
  signal mmio_inst_mmio_rready                              : std_logic;
  signal mmio_inst_mmio_rdata                               : std_logic_vector(31 downto 0);
  signal mmio_inst_mmio_rresp                               : std_logic_vector(1 downto 0);

  signal ss_sold_date_sk_cmd_accm_inst_kernel_cmd_valid     : std_logic;
  signal ss_sold_date_sk_cmd_accm_inst_kernel_cmd_ready     : std_logic;
  signal ss_sold_date_sk_cmd_accm_inst_kernel_cmd_firstIdx  : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal ss_sold_date_sk_cmd_accm_inst_kernel_cmd_lastIdx   : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal ss_sold_date_sk_cmd_accm_inst_kernel_cmd_tag       : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal ss_sold_date_sk_cmd_accm_inst_nucleus_cmd_valid    : std_logic;
  signal ss_sold_date_sk_cmd_accm_inst_nucleus_cmd_ready    : std_logic;
  signal ss_sold_date_sk_cmd_accm_inst_nucleus_cmd_firstIdx : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal ss_sold_date_sk_cmd_accm_inst_nucleus_cmd_lastIdx  : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal ss_sold_date_sk_cmd_accm_inst_nucleus_cmd_ctrl     : std_logic_vector(SS_SOLD_DATE_SK_BUS_ADDR_WIDTH-1 downto 0);
  signal ss_sold_date_sk_cmd_accm_inst_nucleus_cmd_tag      : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal ss_cdemo_sk_cmd_accm_inst_kernel_cmd_valid         : std_logic;
  signal ss_cdemo_sk_cmd_accm_inst_kernel_cmd_ready         : std_logic;
  signal ss_cdemo_sk_cmd_accm_inst_kernel_cmd_firstIdx      : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal ss_cdemo_sk_cmd_accm_inst_kernel_cmd_lastIdx       : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal ss_cdemo_sk_cmd_accm_inst_kernel_cmd_tag           : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal ss_cdemo_sk_cmd_accm_inst_nucleus_cmd_valid        : std_logic;
  signal ss_cdemo_sk_cmd_accm_inst_nucleus_cmd_ready        : std_logic;
  signal ss_cdemo_sk_cmd_accm_inst_nucleus_cmd_firstIdx     : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal ss_cdemo_sk_cmd_accm_inst_nucleus_cmd_lastIdx      : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal ss_cdemo_sk_cmd_accm_inst_nucleus_cmd_ctrl         : std_logic_vector(SS_CDEMO_SK_BUS_ADDR_WIDTH-1 downto 0);
  signal ss_cdemo_sk_cmd_accm_inst_nucleus_cmd_tag          : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal ss_addr_sk_cmd_accm_inst_kernel_cmd_valid          : std_logic;
  signal ss_addr_sk_cmd_accm_inst_kernel_cmd_ready          : std_logic;
  signal ss_addr_sk_cmd_accm_inst_kernel_cmd_firstIdx       : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal ss_addr_sk_cmd_accm_inst_kernel_cmd_lastIdx        : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal ss_addr_sk_cmd_accm_inst_kernel_cmd_tag            : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal ss_addr_sk_cmd_accm_inst_nucleus_cmd_valid         : std_logic;
  signal ss_addr_sk_cmd_accm_inst_nucleus_cmd_ready         : std_logic;
  signal ss_addr_sk_cmd_accm_inst_nucleus_cmd_firstIdx      : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal ss_addr_sk_cmd_accm_inst_nucleus_cmd_lastIdx       : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal ss_addr_sk_cmd_accm_inst_nucleus_cmd_ctrl          : std_logic_vector(SS_ADDR_SK_BUS_ADDR_WIDTH-1 downto 0);
  signal ss_addr_sk_cmd_accm_inst_nucleus_cmd_tag           : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal ss_store_sk_cmd_accm_inst_kernel_cmd_valid         : std_logic;
  signal ss_store_sk_cmd_accm_inst_kernel_cmd_ready         : std_logic;
  signal ss_store_sk_cmd_accm_inst_kernel_cmd_firstIdx      : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal ss_store_sk_cmd_accm_inst_kernel_cmd_lastIdx       : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal ss_store_sk_cmd_accm_inst_kernel_cmd_tag           : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal ss_store_sk_cmd_accm_inst_nucleus_cmd_valid        : std_logic;
  signal ss_store_sk_cmd_accm_inst_nucleus_cmd_ready        : std_logic;
  signal ss_store_sk_cmd_accm_inst_nucleus_cmd_firstIdx     : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal ss_store_sk_cmd_accm_inst_nucleus_cmd_lastIdx      : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal ss_store_sk_cmd_accm_inst_nucleus_cmd_ctrl         : std_logic_vector(SS_STORE_SK_BUS_ADDR_WIDTH-1 downto 0);
  signal ss_store_sk_cmd_accm_inst_nucleus_cmd_tag          : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal ss_quantity_cmd_accm_inst_kernel_cmd_valid         : std_logic;
  signal ss_quantity_cmd_accm_inst_kernel_cmd_ready         : std_logic;
  signal ss_quantity_cmd_accm_inst_kernel_cmd_firstIdx      : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal ss_quantity_cmd_accm_inst_kernel_cmd_lastIdx       : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal ss_quantity_cmd_accm_inst_kernel_cmd_tag           : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal ss_quantity_cmd_accm_inst_nucleus_cmd_valid        : std_logic;
  signal ss_quantity_cmd_accm_inst_nucleus_cmd_ready        : std_logic;
  signal ss_quantity_cmd_accm_inst_nucleus_cmd_firstIdx     : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal ss_quantity_cmd_accm_inst_nucleus_cmd_lastIdx      : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal ss_quantity_cmd_accm_inst_nucleus_cmd_ctrl         : std_logic_vector(SS_QUANTITY_BUS_ADDR_WIDTH-1 downto 0);
  signal ss_quantity_cmd_accm_inst_nucleus_cmd_tag          : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal ss_sales_price_cmd_accm_inst_kernel_cmd_valid      : std_logic;
  signal ss_sales_price_cmd_accm_inst_kernel_cmd_ready      : std_logic;
  signal ss_sales_price_cmd_accm_inst_kernel_cmd_firstIdx   : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal ss_sales_price_cmd_accm_inst_kernel_cmd_lastIdx    : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal ss_sales_price_cmd_accm_inst_kernel_cmd_tag        : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal ss_sales_price_cmd_accm_inst_nucleus_cmd_valid     : std_logic;
  signal ss_sales_price_cmd_accm_inst_nucleus_cmd_ready     : std_logic;
  signal ss_sales_price_cmd_accm_inst_nucleus_cmd_firstIdx  : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal ss_sales_price_cmd_accm_inst_nucleus_cmd_lastIdx   : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal ss_sales_price_cmd_accm_inst_nucleus_cmd_ctrl      : std_logic_vector(SS_SALES_PRICE_BUS_ADDR_WIDTH-1 downto 0);
  signal ss_sales_price_cmd_accm_inst_nucleus_cmd_tag       : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal ss_net_profit_cmd_accm_inst_kernel_cmd_valid       : std_logic;
  signal ss_net_profit_cmd_accm_inst_kernel_cmd_ready       : std_logic;
  signal ss_net_profit_cmd_accm_inst_kernel_cmd_firstIdx    : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal ss_net_profit_cmd_accm_inst_kernel_cmd_lastIdx     : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal ss_net_profit_cmd_accm_inst_kernel_cmd_tag         : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal ss_net_profit_cmd_accm_inst_nucleus_cmd_valid      : std_logic;
  signal ss_net_profit_cmd_accm_inst_nucleus_cmd_ready      : std_logic;
  signal ss_net_profit_cmd_accm_inst_nucleus_cmd_firstIdx   : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal ss_net_profit_cmd_accm_inst_nucleus_cmd_lastIdx    : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal ss_net_profit_cmd_accm_inst_nucleus_cmd_ctrl       : std_logic_vector(SS_NET_PROFIT_BUS_ADDR_WIDTH-1 downto 0);
  signal ss_net_profit_cmd_accm_inst_nucleus_cmd_tag        : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal ss_sold_date_sk_cmd_accm_inst_ctrl : std_logic_vector(SS_SOLD_DATE_SK_BUS_ADDR_WIDTH-1 downto 0);
  signal ss_cdemo_sk_cmd_accm_inst_ctrl     : std_logic_vector(SS_CDEMO_SK_BUS_ADDR_WIDTH-1 downto 0);
  signal ss_addr_sk_cmd_accm_inst_ctrl      : std_logic_vector(SS_ADDR_SK_BUS_ADDR_WIDTH-1 downto 0);
  signal ss_store_sk_cmd_accm_inst_ctrl     : std_logic_vector(SS_STORE_SK_BUS_ADDR_WIDTH-1 downto 0);
  signal ss_quantity_cmd_accm_inst_ctrl     : std_logic_vector(SS_QUANTITY_BUS_ADDR_WIDTH-1 downto 0);
  signal ss_sales_price_cmd_accm_inst_ctrl  : std_logic_vector(SS_SALES_PRICE_BUS_ADDR_WIDTH-1 downto 0);
  signal ss_net_profit_cmd_accm_inst_ctrl   : std_logic_vector(SS_NET_PROFIT_BUS_ADDR_WIDTH-1 downto 0);

begin
  Join_inst : Join
    generic map (
      INDEX_WIDTH => 32,
      TAG_WIDTH   => 1
    )
    port map (
      kcd_clk                      => kcd_clk,
      kcd_reset                    => kcd_reset,
      ss_sold_date_sk_valid        => Join_inst_ss_sold_date_sk_valid,
      ss_sold_date_sk_ready        => Join_inst_ss_sold_date_sk_ready,
      ss_sold_date_sk_dvalid       => Join_inst_ss_sold_date_sk_dvalid,
      ss_sold_date_sk_last         => Join_inst_ss_sold_date_sk_last,
      ss_sold_date_sk              => Join_inst_ss_sold_date_sk,
      ss_cdemo_sk_valid            => Join_inst_ss_cdemo_sk_valid,
      ss_cdemo_sk_ready            => Join_inst_ss_cdemo_sk_ready,
      ss_cdemo_sk_dvalid           => Join_inst_ss_cdemo_sk_dvalid,
      ss_cdemo_sk_last             => Join_inst_ss_cdemo_sk_last,
      ss_cdemo_sk                  => Join_inst_ss_cdemo_sk,
      ss_addr_sk_valid             => Join_inst_ss_addr_sk_valid,
      ss_addr_sk_ready             => Join_inst_ss_addr_sk_ready,
      ss_addr_sk_dvalid            => Join_inst_ss_addr_sk_dvalid,
      ss_addr_sk_last              => Join_inst_ss_addr_sk_last,
      ss_addr_sk                   => Join_inst_ss_addr_sk,
      ss_store_sk_valid            => Join_inst_ss_store_sk_valid,
      ss_store_sk_ready            => Join_inst_ss_store_sk_ready,
      ss_store_sk_dvalid           => Join_inst_ss_store_sk_dvalid,
      ss_store_sk_last             => Join_inst_ss_store_sk_last,
      ss_store_sk                  => Join_inst_ss_store_sk,
      ss_quantity_valid            => Join_inst_ss_quantity_valid,
      ss_quantity_ready            => Join_inst_ss_quantity_ready,
      ss_quantity_dvalid           => Join_inst_ss_quantity_dvalid,
      ss_quantity_last             => Join_inst_ss_quantity_last,
      ss_quantity                  => Join_inst_ss_quantity,
      ss_sales_price_valid         => Join_inst_ss_sales_price_valid,
      ss_sales_price_ready         => Join_inst_ss_sales_price_ready,
      ss_sales_price_dvalid        => Join_inst_ss_sales_price_dvalid,
      ss_sales_price_last          => Join_inst_ss_sales_price_last,
      ss_sales_price               => Join_inst_ss_sales_price,
      ss_net_profit_valid          => Join_inst_ss_net_profit_valid,
      ss_net_profit_ready          => Join_inst_ss_net_profit_ready,
      ss_net_profit_dvalid         => Join_inst_ss_net_profit_dvalid,
      ss_net_profit_last           => Join_inst_ss_net_profit_last,
      ss_net_profit                => Join_inst_ss_net_profit,
      ss_sold_date_sk_unl_valid    => Join_inst_ss_sold_date_sk_unl_valid,
      ss_sold_date_sk_unl_ready    => Join_inst_ss_sold_date_sk_unl_ready,
      ss_sold_date_sk_unl_tag      => Join_inst_ss_sold_date_sk_unl_tag,
      ss_cdemo_sk_unl_valid        => Join_inst_ss_cdemo_sk_unl_valid,
      ss_cdemo_sk_unl_ready        => Join_inst_ss_cdemo_sk_unl_ready,
      ss_cdemo_sk_unl_tag          => Join_inst_ss_cdemo_sk_unl_tag,
      ss_addr_sk_unl_valid         => Join_inst_ss_addr_sk_unl_valid,
      ss_addr_sk_unl_ready         => Join_inst_ss_addr_sk_unl_ready,
      ss_addr_sk_unl_tag           => Join_inst_ss_addr_sk_unl_tag,
      ss_store_sk_unl_valid        => Join_inst_ss_store_sk_unl_valid,
      ss_store_sk_unl_ready        => Join_inst_ss_store_sk_unl_ready,
      ss_store_sk_unl_tag          => Join_inst_ss_store_sk_unl_tag,
      ss_quantity_unl_valid        => Join_inst_ss_quantity_unl_valid,
      ss_quantity_unl_ready        => Join_inst_ss_quantity_unl_ready,
      ss_quantity_unl_tag          => Join_inst_ss_quantity_unl_tag,
      ss_sales_price_unl_valid     => Join_inst_ss_sales_price_unl_valid,
      ss_sales_price_unl_ready     => Join_inst_ss_sales_price_unl_ready,
      ss_sales_price_unl_tag       => Join_inst_ss_sales_price_unl_tag,
      ss_net_profit_unl_valid      => Join_inst_ss_net_profit_unl_valid,
      ss_net_profit_unl_ready      => Join_inst_ss_net_profit_unl_ready,
      ss_net_profit_unl_tag        => Join_inst_ss_net_profit_unl_tag,
      ss_sold_date_sk_cmd_valid    => Join_inst_ss_sold_date_sk_cmd_valid,
      ss_sold_date_sk_cmd_ready    => Join_inst_ss_sold_date_sk_cmd_ready,
      ss_sold_date_sk_cmd_firstIdx => Join_inst_ss_sold_date_sk_cmd_firstIdx,
      ss_sold_date_sk_cmd_lastIdx  => Join_inst_ss_sold_date_sk_cmd_lastIdx,
      ss_sold_date_sk_cmd_tag      => Join_inst_ss_sold_date_sk_cmd_tag,
      ss_cdemo_sk_cmd_valid        => Join_inst_ss_cdemo_sk_cmd_valid,
      ss_cdemo_sk_cmd_ready        => Join_inst_ss_cdemo_sk_cmd_ready,
      ss_cdemo_sk_cmd_firstIdx     => Join_inst_ss_cdemo_sk_cmd_firstIdx,
      ss_cdemo_sk_cmd_lastIdx      => Join_inst_ss_cdemo_sk_cmd_lastIdx,
      ss_cdemo_sk_cmd_tag          => Join_inst_ss_cdemo_sk_cmd_tag,
      ss_addr_sk_cmd_valid         => Join_inst_ss_addr_sk_cmd_valid,
      ss_addr_sk_cmd_ready         => Join_inst_ss_addr_sk_cmd_ready,
      ss_addr_sk_cmd_firstIdx      => Join_inst_ss_addr_sk_cmd_firstIdx,
      ss_addr_sk_cmd_lastIdx       => Join_inst_ss_addr_sk_cmd_lastIdx,
      ss_addr_sk_cmd_tag           => Join_inst_ss_addr_sk_cmd_tag,
      ss_store_sk_cmd_valid        => Join_inst_ss_store_sk_cmd_valid,
      ss_store_sk_cmd_ready        => Join_inst_ss_store_sk_cmd_ready,
      ss_store_sk_cmd_firstIdx     => Join_inst_ss_store_sk_cmd_firstIdx,
      ss_store_sk_cmd_lastIdx      => Join_inst_ss_store_sk_cmd_lastIdx,
      ss_store_sk_cmd_tag          => Join_inst_ss_store_sk_cmd_tag,
      ss_quantity_cmd_valid        => Join_inst_ss_quantity_cmd_valid,
      ss_quantity_cmd_ready        => Join_inst_ss_quantity_cmd_ready,
      ss_quantity_cmd_firstIdx     => Join_inst_ss_quantity_cmd_firstIdx,
      ss_quantity_cmd_lastIdx      => Join_inst_ss_quantity_cmd_lastIdx,
      ss_quantity_cmd_tag          => Join_inst_ss_quantity_cmd_tag,
      ss_sales_price_cmd_valid     => Join_inst_ss_sales_price_cmd_valid,
      ss_sales_price_cmd_ready     => Join_inst_ss_sales_price_cmd_ready,
      ss_sales_price_cmd_firstIdx  => Join_inst_ss_sales_price_cmd_firstIdx,
      ss_sales_price_cmd_lastIdx   => Join_inst_ss_sales_price_cmd_lastIdx,
      ss_sales_price_cmd_tag       => Join_inst_ss_sales_price_cmd_tag,
      ss_net_profit_cmd_valid      => Join_inst_ss_net_profit_cmd_valid,
      ss_net_profit_cmd_ready      => Join_inst_ss_net_profit_cmd_ready,
      ss_net_profit_cmd_firstIdx   => Join_inst_ss_net_profit_cmd_firstIdx,
      ss_net_profit_cmd_lastIdx    => Join_inst_ss_net_profit_cmd_lastIdx,
      ss_net_profit_cmd_tag        => Join_inst_ss_net_profit_cmd_tag,
      start                        => Join_inst_start,
      stop                         => Join_inst_stop,
      reset                        => Join_inst_reset,
      idle                         => Join_inst_idle,
      busy                         => Join_inst_busy,
      done                         => Join_inst_done,
      result                       => Join_inst_result,
      ss_firstidx                  => Join_inst_ss_firstidx,
      ss_lastidx                   => Join_inst_ss_lastidx
    );

  mmio_inst : mmio
    port map (
      kcd_clk                       => kcd_clk,
      kcd_reset                     => kcd_reset,
      f_start_data                  => mmio_inst_f_start_data,
      f_stop_data                   => mmio_inst_f_stop_data,
      f_reset_data                  => mmio_inst_f_reset_data,
      f_idle_write_data             => mmio_inst_f_idle_write_data,
      f_busy_write_data             => mmio_inst_f_busy_write_data,
      f_done_write_data             => mmio_inst_f_done_write_data,
      f_result_write_data           => mmio_inst_f_result_write_data,
      f_ss_firstidx_data            => mmio_inst_f_ss_firstidx_data,
      f_ss_lastidx_data             => mmio_inst_f_ss_lastidx_data,
      f_ss_sold_date_sk_values_data => mmio_inst_f_ss_sold_date_sk_values_data,
      f_ss_cdemo_sk_values_data     => mmio_inst_f_ss_cdemo_sk_values_data,
      f_ss_addr_sk_values_data      => mmio_inst_f_ss_addr_sk_values_data,
      f_ss_store_sk_values_data     => mmio_inst_f_ss_store_sk_values_data,
      f_ss_quantity_values_data     => mmio_inst_f_ss_quantity_values_data,
      f_ss_sales_price_values_data  => mmio_inst_f_ss_sales_price_values_data,
      f_ss_net_profit_values_data   => mmio_inst_f_ss_net_profit_values_data,
      mmio_awvalid                  => mmio_inst_mmio_awvalid,
      mmio_awready                  => mmio_inst_mmio_awready,
      mmio_awaddr                   => mmio_inst_mmio_awaddr,
      mmio_wvalid                   => mmio_inst_mmio_wvalid,
      mmio_wready                   => mmio_inst_mmio_wready,
      mmio_wdata                    => mmio_inst_mmio_wdata,
      mmio_wstrb                    => mmio_inst_mmio_wstrb,
      mmio_bvalid                   => mmio_inst_mmio_bvalid,
      mmio_bready                   => mmio_inst_mmio_bready,
      mmio_bresp                    => mmio_inst_mmio_bresp,
      mmio_arvalid                  => mmio_inst_mmio_arvalid,
      mmio_arready                  => mmio_inst_mmio_arready,
      mmio_araddr                   => mmio_inst_mmio_araddr,
      mmio_rvalid                   => mmio_inst_mmio_rvalid,
      mmio_rready                   => mmio_inst_mmio_rready,
      mmio_rdata                    => mmio_inst_mmio_rdata,
      mmio_rresp                    => mmio_inst_mmio_rresp
    );

  ss_sold_date_sk_cmd_accm_inst : ArrayCmdCtrlMerger
    generic map (
      NUM_ADDR       => 1,
      BUS_ADDR_WIDTH => SS_SOLD_DATE_SK_BUS_ADDR_WIDTH,
      INDEX_WIDTH    => INDEX_WIDTH,
      TAG_WIDTH      => TAG_WIDTH
    )
    port map (
      kernel_cmd_valid     => ss_sold_date_sk_cmd_accm_inst_kernel_cmd_valid,
      kernel_cmd_ready     => ss_sold_date_sk_cmd_accm_inst_kernel_cmd_ready,
      kernel_cmd_firstIdx  => ss_sold_date_sk_cmd_accm_inst_kernel_cmd_firstIdx,
      kernel_cmd_lastIdx   => ss_sold_date_sk_cmd_accm_inst_kernel_cmd_lastIdx,
      kernel_cmd_tag       => ss_sold_date_sk_cmd_accm_inst_kernel_cmd_tag,
      nucleus_cmd_valid    => ss_sold_date_sk_cmd_accm_inst_nucleus_cmd_valid,
      nucleus_cmd_ready    => ss_sold_date_sk_cmd_accm_inst_nucleus_cmd_ready,
      nucleus_cmd_firstIdx => ss_sold_date_sk_cmd_accm_inst_nucleus_cmd_firstIdx,
      nucleus_cmd_lastIdx  => ss_sold_date_sk_cmd_accm_inst_nucleus_cmd_lastIdx,
      nucleus_cmd_ctrl     => ss_sold_date_sk_cmd_accm_inst_nucleus_cmd_ctrl,
      nucleus_cmd_tag      => ss_sold_date_sk_cmd_accm_inst_nucleus_cmd_tag,
      ctrl                 => ss_sold_date_sk_cmd_accm_inst_ctrl
    );

  ss_cdemo_sk_cmd_accm_inst : ArrayCmdCtrlMerger
    generic map (
      NUM_ADDR       => 1,
      BUS_ADDR_WIDTH => SS_CDEMO_SK_BUS_ADDR_WIDTH,
      INDEX_WIDTH    => INDEX_WIDTH,
      TAG_WIDTH      => TAG_WIDTH
    )
    port map (
      kernel_cmd_valid     => ss_cdemo_sk_cmd_accm_inst_kernel_cmd_valid,
      kernel_cmd_ready     => ss_cdemo_sk_cmd_accm_inst_kernel_cmd_ready,
      kernel_cmd_firstIdx  => ss_cdemo_sk_cmd_accm_inst_kernel_cmd_firstIdx,
      kernel_cmd_lastIdx   => ss_cdemo_sk_cmd_accm_inst_kernel_cmd_lastIdx,
      kernel_cmd_tag       => ss_cdemo_sk_cmd_accm_inst_kernel_cmd_tag,
      nucleus_cmd_valid    => ss_cdemo_sk_cmd_accm_inst_nucleus_cmd_valid,
      nucleus_cmd_ready    => ss_cdemo_sk_cmd_accm_inst_nucleus_cmd_ready,
      nucleus_cmd_firstIdx => ss_cdemo_sk_cmd_accm_inst_nucleus_cmd_firstIdx,
      nucleus_cmd_lastIdx  => ss_cdemo_sk_cmd_accm_inst_nucleus_cmd_lastIdx,
      nucleus_cmd_ctrl     => ss_cdemo_sk_cmd_accm_inst_nucleus_cmd_ctrl,
      nucleus_cmd_tag      => ss_cdemo_sk_cmd_accm_inst_nucleus_cmd_tag,
      ctrl                 => ss_cdemo_sk_cmd_accm_inst_ctrl
    );

  ss_addr_sk_cmd_accm_inst : ArrayCmdCtrlMerger
    generic map (
      NUM_ADDR       => 1,
      BUS_ADDR_WIDTH => SS_ADDR_SK_BUS_ADDR_WIDTH,
      INDEX_WIDTH    => INDEX_WIDTH,
      TAG_WIDTH      => TAG_WIDTH
    )
    port map (
      kernel_cmd_valid     => ss_addr_sk_cmd_accm_inst_kernel_cmd_valid,
      kernel_cmd_ready     => ss_addr_sk_cmd_accm_inst_kernel_cmd_ready,
      kernel_cmd_firstIdx  => ss_addr_sk_cmd_accm_inst_kernel_cmd_firstIdx,
      kernel_cmd_lastIdx   => ss_addr_sk_cmd_accm_inst_kernel_cmd_lastIdx,
      kernel_cmd_tag       => ss_addr_sk_cmd_accm_inst_kernel_cmd_tag,
      nucleus_cmd_valid    => ss_addr_sk_cmd_accm_inst_nucleus_cmd_valid,
      nucleus_cmd_ready    => ss_addr_sk_cmd_accm_inst_nucleus_cmd_ready,
      nucleus_cmd_firstIdx => ss_addr_sk_cmd_accm_inst_nucleus_cmd_firstIdx,
      nucleus_cmd_lastIdx  => ss_addr_sk_cmd_accm_inst_nucleus_cmd_lastIdx,
      nucleus_cmd_ctrl     => ss_addr_sk_cmd_accm_inst_nucleus_cmd_ctrl,
      nucleus_cmd_tag      => ss_addr_sk_cmd_accm_inst_nucleus_cmd_tag,
      ctrl                 => ss_addr_sk_cmd_accm_inst_ctrl
    );

  ss_store_sk_cmd_accm_inst : ArrayCmdCtrlMerger
    generic map (
      NUM_ADDR       => 1,
      BUS_ADDR_WIDTH => SS_STORE_SK_BUS_ADDR_WIDTH,
      INDEX_WIDTH    => INDEX_WIDTH,
      TAG_WIDTH      => TAG_WIDTH
    )
    port map (
      kernel_cmd_valid     => ss_store_sk_cmd_accm_inst_kernel_cmd_valid,
      kernel_cmd_ready     => ss_store_sk_cmd_accm_inst_kernel_cmd_ready,
      kernel_cmd_firstIdx  => ss_store_sk_cmd_accm_inst_kernel_cmd_firstIdx,
      kernel_cmd_lastIdx   => ss_store_sk_cmd_accm_inst_kernel_cmd_lastIdx,
      kernel_cmd_tag       => ss_store_sk_cmd_accm_inst_kernel_cmd_tag,
      nucleus_cmd_valid    => ss_store_sk_cmd_accm_inst_nucleus_cmd_valid,
      nucleus_cmd_ready    => ss_store_sk_cmd_accm_inst_nucleus_cmd_ready,
      nucleus_cmd_firstIdx => ss_store_sk_cmd_accm_inst_nucleus_cmd_firstIdx,
      nucleus_cmd_lastIdx  => ss_store_sk_cmd_accm_inst_nucleus_cmd_lastIdx,
      nucleus_cmd_ctrl     => ss_store_sk_cmd_accm_inst_nucleus_cmd_ctrl,
      nucleus_cmd_tag      => ss_store_sk_cmd_accm_inst_nucleus_cmd_tag,
      ctrl                 => ss_store_sk_cmd_accm_inst_ctrl
    );

  ss_quantity_cmd_accm_inst : ArrayCmdCtrlMerger
    generic map (
      NUM_ADDR       => 1,
      BUS_ADDR_WIDTH => SS_QUANTITY_BUS_ADDR_WIDTH,
      INDEX_WIDTH    => INDEX_WIDTH,
      TAG_WIDTH      => TAG_WIDTH
    )
    port map (
      kernel_cmd_valid     => ss_quantity_cmd_accm_inst_kernel_cmd_valid,
      kernel_cmd_ready     => ss_quantity_cmd_accm_inst_kernel_cmd_ready,
      kernel_cmd_firstIdx  => ss_quantity_cmd_accm_inst_kernel_cmd_firstIdx,
      kernel_cmd_lastIdx   => ss_quantity_cmd_accm_inst_kernel_cmd_lastIdx,
      kernel_cmd_tag       => ss_quantity_cmd_accm_inst_kernel_cmd_tag,
      nucleus_cmd_valid    => ss_quantity_cmd_accm_inst_nucleus_cmd_valid,
      nucleus_cmd_ready    => ss_quantity_cmd_accm_inst_nucleus_cmd_ready,
      nucleus_cmd_firstIdx => ss_quantity_cmd_accm_inst_nucleus_cmd_firstIdx,
      nucleus_cmd_lastIdx  => ss_quantity_cmd_accm_inst_nucleus_cmd_lastIdx,
      nucleus_cmd_ctrl     => ss_quantity_cmd_accm_inst_nucleus_cmd_ctrl,
      nucleus_cmd_tag      => ss_quantity_cmd_accm_inst_nucleus_cmd_tag,
      ctrl                 => ss_quantity_cmd_accm_inst_ctrl
    );

  ss_sales_price_cmd_accm_inst : ArrayCmdCtrlMerger
    generic map (
      NUM_ADDR       => 1,
      BUS_ADDR_WIDTH => SS_SALES_PRICE_BUS_ADDR_WIDTH,
      INDEX_WIDTH    => INDEX_WIDTH,
      TAG_WIDTH      => TAG_WIDTH
    )
    port map (
      kernel_cmd_valid     => ss_sales_price_cmd_accm_inst_kernel_cmd_valid,
      kernel_cmd_ready     => ss_sales_price_cmd_accm_inst_kernel_cmd_ready,
      kernel_cmd_firstIdx  => ss_sales_price_cmd_accm_inst_kernel_cmd_firstIdx,
      kernel_cmd_lastIdx   => ss_sales_price_cmd_accm_inst_kernel_cmd_lastIdx,
      kernel_cmd_tag       => ss_sales_price_cmd_accm_inst_kernel_cmd_tag,
      nucleus_cmd_valid    => ss_sales_price_cmd_accm_inst_nucleus_cmd_valid,
      nucleus_cmd_ready    => ss_sales_price_cmd_accm_inst_nucleus_cmd_ready,
      nucleus_cmd_firstIdx => ss_sales_price_cmd_accm_inst_nucleus_cmd_firstIdx,
      nucleus_cmd_lastIdx  => ss_sales_price_cmd_accm_inst_nucleus_cmd_lastIdx,
      nucleus_cmd_ctrl     => ss_sales_price_cmd_accm_inst_nucleus_cmd_ctrl,
      nucleus_cmd_tag      => ss_sales_price_cmd_accm_inst_nucleus_cmd_tag,
      ctrl                 => ss_sales_price_cmd_accm_inst_ctrl
    );

  ss_net_profit_cmd_accm_inst : ArrayCmdCtrlMerger
    generic map (
      NUM_ADDR       => 1,
      BUS_ADDR_WIDTH => SS_NET_PROFIT_BUS_ADDR_WIDTH,
      INDEX_WIDTH    => INDEX_WIDTH,
      TAG_WIDTH      => TAG_WIDTH
    )
    port map (
      kernel_cmd_valid     => ss_net_profit_cmd_accm_inst_kernel_cmd_valid,
      kernel_cmd_ready     => ss_net_profit_cmd_accm_inst_kernel_cmd_ready,
      kernel_cmd_firstIdx  => ss_net_profit_cmd_accm_inst_kernel_cmd_firstIdx,
      kernel_cmd_lastIdx   => ss_net_profit_cmd_accm_inst_kernel_cmd_lastIdx,
      kernel_cmd_tag       => ss_net_profit_cmd_accm_inst_kernel_cmd_tag,
      nucleus_cmd_valid    => ss_net_profit_cmd_accm_inst_nucleus_cmd_valid,
      nucleus_cmd_ready    => ss_net_profit_cmd_accm_inst_nucleus_cmd_ready,
      nucleus_cmd_firstIdx => ss_net_profit_cmd_accm_inst_nucleus_cmd_firstIdx,
      nucleus_cmd_lastIdx  => ss_net_profit_cmd_accm_inst_nucleus_cmd_lastIdx,
      nucleus_cmd_ctrl     => ss_net_profit_cmd_accm_inst_nucleus_cmd_ctrl,
      nucleus_cmd_tag      => ss_net_profit_cmd_accm_inst_nucleus_cmd_tag,
      ctrl                 => ss_net_profit_cmd_accm_inst_ctrl
    );

  ss_sold_date_sk_cmd_valid                       <= ss_sold_date_sk_cmd_accm_inst_nucleus_cmd_valid;
  ss_sold_date_sk_cmd_accm_inst_nucleus_cmd_ready <= ss_sold_date_sk_cmd_ready;
  ss_sold_date_sk_cmd_firstIdx                    <= ss_sold_date_sk_cmd_accm_inst_nucleus_cmd_firstIdx;
  ss_sold_date_sk_cmd_lastIdx                     <= ss_sold_date_sk_cmd_accm_inst_nucleus_cmd_lastIdx;
  ss_sold_date_sk_cmd_ctrl                        <= ss_sold_date_sk_cmd_accm_inst_nucleus_cmd_ctrl;
  ss_sold_date_sk_cmd_tag                         <= ss_sold_date_sk_cmd_accm_inst_nucleus_cmd_tag;

  ss_cdemo_sk_cmd_valid                           <= ss_cdemo_sk_cmd_accm_inst_nucleus_cmd_valid;
  ss_cdemo_sk_cmd_accm_inst_nucleus_cmd_ready     <= ss_cdemo_sk_cmd_ready;
  ss_cdemo_sk_cmd_firstIdx                        <= ss_cdemo_sk_cmd_accm_inst_nucleus_cmd_firstIdx;
  ss_cdemo_sk_cmd_lastIdx                         <= ss_cdemo_sk_cmd_accm_inst_nucleus_cmd_lastIdx;
  ss_cdemo_sk_cmd_ctrl                            <= ss_cdemo_sk_cmd_accm_inst_nucleus_cmd_ctrl;
  ss_cdemo_sk_cmd_tag                             <= ss_cdemo_sk_cmd_accm_inst_nucleus_cmd_tag;

  ss_addr_sk_cmd_valid                            <= ss_addr_sk_cmd_accm_inst_nucleus_cmd_valid;
  ss_addr_sk_cmd_accm_inst_nucleus_cmd_ready      <= ss_addr_sk_cmd_ready;
  ss_addr_sk_cmd_firstIdx                         <= ss_addr_sk_cmd_accm_inst_nucleus_cmd_firstIdx;
  ss_addr_sk_cmd_lastIdx                          <= ss_addr_sk_cmd_accm_inst_nucleus_cmd_lastIdx;
  ss_addr_sk_cmd_ctrl                             <= ss_addr_sk_cmd_accm_inst_nucleus_cmd_ctrl;
  ss_addr_sk_cmd_tag                              <= ss_addr_sk_cmd_accm_inst_nucleus_cmd_tag;

  ss_store_sk_cmd_valid                           <= ss_store_sk_cmd_accm_inst_nucleus_cmd_valid;
  ss_store_sk_cmd_accm_inst_nucleus_cmd_ready     <= ss_store_sk_cmd_ready;
  ss_store_sk_cmd_firstIdx                        <= ss_store_sk_cmd_accm_inst_nucleus_cmd_firstIdx;
  ss_store_sk_cmd_lastIdx                         <= ss_store_sk_cmd_accm_inst_nucleus_cmd_lastIdx;
  ss_store_sk_cmd_ctrl                            <= ss_store_sk_cmd_accm_inst_nucleus_cmd_ctrl;
  ss_store_sk_cmd_tag                             <= ss_store_sk_cmd_accm_inst_nucleus_cmd_tag;

  ss_quantity_cmd_valid                           <= ss_quantity_cmd_accm_inst_nucleus_cmd_valid;
  ss_quantity_cmd_accm_inst_nucleus_cmd_ready     <= ss_quantity_cmd_ready;
  ss_quantity_cmd_firstIdx                        <= ss_quantity_cmd_accm_inst_nucleus_cmd_firstIdx;
  ss_quantity_cmd_lastIdx                         <= ss_quantity_cmd_accm_inst_nucleus_cmd_lastIdx;
  ss_quantity_cmd_ctrl                            <= ss_quantity_cmd_accm_inst_nucleus_cmd_ctrl;
  ss_quantity_cmd_tag                             <= ss_quantity_cmd_accm_inst_nucleus_cmd_tag;

  ss_sales_price_cmd_valid                        <= ss_sales_price_cmd_accm_inst_nucleus_cmd_valid;
  ss_sales_price_cmd_accm_inst_nucleus_cmd_ready  <= ss_sales_price_cmd_ready;
  ss_sales_price_cmd_firstIdx                     <= ss_sales_price_cmd_accm_inst_nucleus_cmd_firstIdx;
  ss_sales_price_cmd_lastIdx                      <= ss_sales_price_cmd_accm_inst_nucleus_cmd_lastIdx;
  ss_sales_price_cmd_ctrl                         <= ss_sales_price_cmd_accm_inst_nucleus_cmd_ctrl;
  ss_sales_price_cmd_tag                          <= ss_sales_price_cmd_accm_inst_nucleus_cmd_tag;

  ss_net_profit_cmd_valid                         <= ss_net_profit_cmd_accm_inst_nucleus_cmd_valid;
  ss_net_profit_cmd_accm_inst_nucleus_cmd_ready   <= ss_net_profit_cmd_ready;
  ss_net_profit_cmd_firstIdx                      <= ss_net_profit_cmd_accm_inst_nucleus_cmd_firstIdx;
  ss_net_profit_cmd_lastIdx                       <= ss_net_profit_cmd_accm_inst_nucleus_cmd_lastIdx;
  ss_net_profit_cmd_ctrl                          <= ss_net_profit_cmd_accm_inst_nucleus_cmd_ctrl;
  ss_net_profit_cmd_tag                           <= ss_net_profit_cmd_accm_inst_nucleus_cmd_tag;

  Join_inst_ss_sold_date_sk_valid                   <= ss_sold_date_sk_valid;
  ss_sold_date_sk_ready                             <= Join_inst_ss_sold_date_sk_ready;
  Join_inst_ss_sold_date_sk_dvalid                  <= ss_sold_date_sk_dvalid;
  Join_inst_ss_sold_date_sk_last                    <= ss_sold_date_sk_last;
  Join_inst_ss_sold_date_sk                         <= ss_sold_date_sk;

  Join_inst_ss_cdemo_sk_valid                       <= ss_cdemo_sk_valid;
  ss_cdemo_sk_ready                                 <= Join_inst_ss_cdemo_sk_ready;
  Join_inst_ss_cdemo_sk_dvalid                      <= ss_cdemo_sk_dvalid;
  Join_inst_ss_cdemo_sk_last                        <= ss_cdemo_sk_last;
  Join_inst_ss_cdemo_sk                             <= ss_cdemo_sk;

  Join_inst_ss_addr_sk_valid                        <= ss_addr_sk_valid;
  ss_addr_sk_ready                                  <= Join_inst_ss_addr_sk_ready;
  Join_inst_ss_addr_sk_dvalid                       <= ss_addr_sk_dvalid;
  Join_inst_ss_addr_sk_last                         <= ss_addr_sk_last;
  Join_inst_ss_addr_sk                              <= ss_addr_sk;

  Join_inst_ss_store_sk_valid                       <= ss_store_sk_valid;
  ss_store_sk_ready                                 <= Join_inst_ss_store_sk_ready;
  Join_inst_ss_store_sk_dvalid                      <= ss_store_sk_dvalid;
  Join_inst_ss_store_sk_last                        <= ss_store_sk_last;
  Join_inst_ss_store_sk                             <= ss_store_sk;

  Join_inst_ss_quantity_valid                       <= ss_quantity_valid;
  ss_quantity_ready                                 <= Join_inst_ss_quantity_ready;
  Join_inst_ss_quantity_dvalid                      <= ss_quantity_dvalid;
  Join_inst_ss_quantity_last                        <= ss_quantity_last;
  Join_inst_ss_quantity                             <= ss_quantity;

  Join_inst_ss_sales_price_valid                    <= ss_sales_price_valid;
  ss_sales_price_ready                              <= Join_inst_ss_sales_price_ready;
  Join_inst_ss_sales_price_dvalid                   <= ss_sales_price_dvalid;
  Join_inst_ss_sales_price_last                     <= ss_sales_price_last;
  Join_inst_ss_sales_price                          <= ss_sales_price;

  Join_inst_ss_net_profit_valid                     <= ss_net_profit_valid;
  ss_net_profit_ready                               <= Join_inst_ss_net_profit_ready;
  Join_inst_ss_net_profit_dvalid                    <= ss_net_profit_dvalid;
  Join_inst_ss_net_profit_last                      <= ss_net_profit_last;
  Join_inst_ss_net_profit                           <= ss_net_profit;

  Join_inst_ss_sold_date_sk_unl_valid               <= ss_sold_date_sk_unl_valid;
  ss_sold_date_sk_unl_ready                         <= Join_inst_ss_sold_date_sk_unl_ready;
  Join_inst_ss_sold_date_sk_unl_tag                 <= ss_sold_date_sk_unl_tag;

  Join_inst_ss_cdemo_sk_unl_valid                   <= ss_cdemo_sk_unl_valid;
  ss_cdemo_sk_unl_ready                             <= Join_inst_ss_cdemo_sk_unl_ready;
  Join_inst_ss_cdemo_sk_unl_tag                     <= ss_cdemo_sk_unl_tag;

  Join_inst_ss_addr_sk_unl_valid                    <= ss_addr_sk_unl_valid;
  ss_addr_sk_unl_ready                              <= Join_inst_ss_addr_sk_unl_ready;
  Join_inst_ss_addr_sk_unl_tag                      <= ss_addr_sk_unl_tag;

  Join_inst_ss_store_sk_unl_valid                   <= ss_store_sk_unl_valid;
  ss_store_sk_unl_ready                             <= Join_inst_ss_store_sk_unl_ready;
  Join_inst_ss_store_sk_unl_tag                     <= ss_store_sk_unl_tag;

  Join_inst_ss_quantity_unl_valid                   <= ss_quantity_unl_valid;
  ss_quantity_unl_ready                             <= Join_inst_ss_quantity_unl_ready;
  Join_inst_ss_quantity_unl_tag                     <= ss_quantity_unl_tag;

  Join_inst_ss_sales_price_unl_valid                <= ss_sales_price_unl_valid;
  ss_sales_price_unl_ready                          <= Join_inst_ss_sales_price_unl_ready;
  Join_inst_ss_sales_price_unl_tag                  <= ss_sales_price_unl_tag;

  Join_inst_ss_net_profit_unl_valid                 <= ss_net_profit_unl_valid;
  ss_net_profit_unl_ready                           <= Join_inst_ss_net_profit_unl_ready;
  Join_inst_ss_net_profit_unl_tag                   <= ss_net_profit_unl_tag;

  Join_inst_start                                   <= mmio_inst_f_start_data;
  Join_inst_stop                                    <= mmio_inst_f_stop_data;
  Join_inst_reset                                   <= mmio_inst_f_reset_data;
  Join_inst_ss_firstidx                             <= mmio_inst_f_ss_firstidx_data;
  Join_inst_ss_lastidx                              <= mmio_inst_f_ss_lastidx_data;
  mmio_inst_f_idle_write_data                       <= Join_inst_idle;
  mmio_inst_f_busy_write_data                       <= Join_inst_busy;
  mmio_inst_f_done_write_data                       <= Join_inst_done;
  mmio_inst_f_result_write_data                     <= Join_inst_result;
  mmio_inst_mmio_awvalid                            <= mmio_awvalid;
  mmio_awready                                      <= mmio_inst_mmio_awready;
  mmio_inst_mmio_awaddr                             <= mmio_awaddr;
  mmio_inst_mmio_wvalid                             <= mmio_wvalid;
  mmio_wready                                       <= mmio_inst_mmio_wready;
  mmio_inst_mmio_wdata                              <= mmio_wdata;
  mmio_inst_mmio_wstrb                              <= mmio_wstrb;
  mmio_bvalid                                       <= mmio_inst_mmio_bvalid;
  mmio_inst_mmio_bready                             <= mmio_bready;
  mmio_bresp                                        <= mmio_inst_mmio_bresp;
  mmio_inst_mmio_arvalid                            <= mmio_arvalid;
  mmio_arready                                      <= mmio_inst_mmio_arready;
  mmio_inst_mmio_araddr                             <= mmio_araddr;
  mmio_rvalid                                       <= mmio_inst_mmio_rvalid;
  mmio_inst_mmio_rready                             <= mmio_rready;
  mmio_rdata                                        <= mmio_inst_mmio_rdata;
  mmio_rresp                                        <= mmio_inst_mmio_rresp;

  ss_sold_date_sk_cmd_accm_inst_kernel_cmd_valid    <= Join_inst_ss_sold_date_sk_cmd_valid;
  Join_inst_ss_sold_date_sk_cmd_ready               <= ss_sold_date_sk_cmd_accm_inst_kernel_cmd_ready;
  ss_sold_date_sk_cmd_accm_inst_kernel_cmd_firstIdx <= Join_inst_ss_sold_date_sk_cmd_firstIdx;
  ss_sold_date_sk_cmd_accm_inst_kernel_cmd_lastIdx  <= Join_inst_ss_sold_date_sk_cmd_lastIdx;
  ss_sold_date_sk_cmd_accm_inst_kernel_cmd_tag      <= Join_inst_ss_sold_date_sk_cmd_tag;

  ss_cdemo_sk_cmd_accm_inst_kernel_cmd_valid        <= Join_inst_ss_cdemo_sk_cmd_valid;
  Join_inst_ss_cdemo_sk_cmd_ready                   <= ss_cdemo_sk_cmd_accm_inst_kernel_cmd_ready;
  ss_cdemo_sk_cmd_accm_inst_kernel_cmd_firstIdx     <= Join_inst_ss_cdemo_sk_cmd_firstIdx;
  ss_cdemo_sk_cmd_accm_inst_kernel_cmd_lastIdx      <= Join_inst_ss_cdemo_sk_cmd_lastIdx;
  ss_cdemo_sk_cmd_accm_inst_kernel_cmd_tag          <= Join_inst_ss_cdemo_sk_cmd_tag;

  ss_addr_sk_cmd_accm_inst_kernel_cmd_valid         <= Join_inst_ss_addr_sk_cmd_valid;
  Join_inst_ss_addr_sk_cmd_ready                    <= ss_addr_sk_cmd_accm_inst_kernel_cmd_ready;
  ss_addr_sk_cmd_accm_inst_kernel_cmd_firstIdx      <= Join_inst_ss_addr_sk_cmd_firstIdx;
  ss_addr_sk_cmd_accm_inst_kernel_cmd_lastIdx       <= Join_inst_ss_addr_sk_cmd_lastIdx;
  ss_addr_sk_cmd_accm_inst_kernel_cmd_tag           <= Join_inst_ss_addr_sk_cmd_tag;

  ss_store_sk_cmd_accm_inst_kernel_cmd_valid        <= Join_inst_ss_store_sk_cmd_valid;
  Join_inst_ss_store_sk_cmd_ready                   <= ss_store_sk_cmd_accm_inst_kernel_cmd_ready;
  ss_store_sk_cmd_accm_inst_kernel_cmd_firstIdx     <= Join_inst_ss_store_sk_cmd_firstIdx;
  ss_store_sk_cmd_accm_inst_kernel_cmd_lastIdx      <= Join_inst_ss_store_sk_cmd_lastIdx;
  ss_store_sk_cmd_accm_inst_kernel_cmd_tag          <= Join_inst_ss_store_sk_cmd_tag;

  ss_quantity_cmd_accm_inst_kernel_cmd_valid        <= Join_inst_ss_quantity_cmd_valid;
  Join_inst_ss_quantity_cmd_ready                   <= ss_quantity_cmd_accm_inst_kernel_cmd_ready;
  ss_quantity_cmd_accm_inst_kernel_cmd_firstIdx     <= Join_inst_ss_quantity_cmd_firstIdx;
  ss_quantity_cmd_accm_inst_kernel_cmd_lastIdx      <= Join_inst_ss_quantity_cmd_lastIdx;
  ss_quantity_cmd_accm_inst_kernel_cmd_tag          <= Join_inst_ss_quantity_cmd_tag;

  ss_sales_price_cmd_accm_inst_kernel_cmd_valid     <= Join_inst_ss_sales_price_cmd_valid;
  Join_inst_ss_sales_price_cmd_ready                <= ss_sales_price_cmd_accm_inst_kernel_cmd_ready;
  ss_sales_price_cmd_accm_inst_kernel_cmd_firstIdx  <= Join_inst_ss_sales_price_cmd_firstIdx;
  ss_sales_price_cmd_accm_inst_kernel_cmd_lastIdx   <= Join_inst_ss_sales_price_cmd_lastIdx;
  ss_sales_price_cmd_accm_inst_kernel_cmd_tag       <= Join_inst_ss_sales_price_cmd_tag;

  ss_net_profit_cmd_accm_inst_kernel_cmd_valid      <= Join_inst_ss_net_profit_cmd_valid;
  Join_inst_ss_net_profit_cmd_ready                 <= ss_net_profit_cmd_accm_inst_kernel_cmd_ready;
  ss_net_profit_cmd_accm_inst_kernel_cmd_firstIdx   <= Join_inst_ss_net_profit_cmd_firstIdx;
  ss_net_profit_cmd_accm_inst_kernel_cmd_lastIdx    <= Join_inst_ss_net_profit_cmd_lastIdx;
  ss_net_profit_cmd_accm_inst_kernel_cmd_tag        <= Join_inst_ss_net_profit_cmd_tag;

  ss_sold_date_sk_cmd_accm_inst_ctrl(63 downto 0) <= mmio_inst_f_ss_sold_date_sk_values_data;
  ss_cdemo_sk_cmd_accm_inst_ctrl(63 downto 0)     <= mmio_inst_f_ss_cdemo_sk_values_data;
  ss_addr_sk_cmd_accm_inst_ctrl(63 downto 0)      <= mmio_inst_f_ss_addr_sk_values_data;
  ss_store_sk_cmd_accm_inst_ctrl(63 downto 0)     <= mmio_inst_f_ss_store_sk_values_data;
  ss_quantity_cmd_accm_inst_ctrl(63 downto 0)     <= mmio_inst_f_ss_quantity_values_data;
  ss_sales_price_cmd_accm_inst_ctrl(63 downto 0)  <= mmio_inst_f_ss_sales_price_values_data;
  ss_net_profit_cmd_accm_inst_ctrl(63 downto 0)   <= mmio_inst_f_ss_net_profit_values_data;

end architecture;
