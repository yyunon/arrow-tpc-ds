-- Copyright 2018-2019 Delft University of Technology
--
-- Licensed under the Apache License, Version 2.0 (the "License");
-- you may not use this file except in compliance with the License.
-- You may obtain a copy of the License at
--
--     http://www.apache.org/licenses/LICENSE-2.0
--
-- Unless required by applicable law or agreed to in writing, software
-- distributed under the License is distributed on an "AS IS" BASIS,
-- WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
-- See the License for the specific language governing permissions and
-- limitations under the License.
--
-- This file was generated by Fletchgen. Modify this file at your own risk.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library work;
use work.Interconnect_pkg.all;

entity Join_Mantle is
  generic (
    INDEX_WIDTH        : integer := 32;
    TAG_WIDTH          : integer := 1;
    BUS_ADDR_WIDTH     : integer := 64;
    BUS_DATA_WIDTH     : integer := 512;
    BUS_LEN_WIDTH      : integer := 8;
    BUS_BURST_STEP_LEN : integer := 1;
    BUS_BURST_MAX_LEN  : integer := 16
  );
  port (
    bcd_clk           : in  std_logic;
    bcd_reset         : in  std_logic;
    kcd_clk           : in  std_logic;
    kcd_reset         : in  std_logic;
    mmio_awvalid      : in  std_logic;
    mmio_awready      : out std_logic;
    mmio_awaddr       : in  std_logic_vector(31 downto 0);
    mmio_wvalid       : in  std_logic;
    mmio_wready       : out std_logic;
    mmio_wdata        : in  std_logic_vector(31 downto 0);
    mmio_wstrb        : in  std_logic_vector(3 downto 0);
    mmio_bvalid       : out std_logic;
    mmio_bready       : in  std_logic;
    mmio_bresp        : out std_logic_vector(1 downto 0);
    mmio_arvalid      : in  std_logic;
    mmio_arready      : out std_logic;
    mmio_araddr       : in  std_logic_vector(31 downto 0);
    mmio_rvalid       : out std_logic;
    mmio_rready       : in  std_logic;
    mmio_rdata        : out std_logic_vector(31 downto 0);
    mmio_rresp        : out std_logic_vector(1 downto 0);
    rd_mst_rreq_valid : out std_logic;
    rd_mst_rreq_ready : in  std_logic;
    rd_mst_rreq_addr  : out std_logic_vector(BUS_ADDR_WIDTH-1 downto 0);
    rd_mst_rreq_len   : out std_logic_vector(BUS_LEN_WIDTH-1 downto 0);
    rd_mst_rdat_valid : in  std_logic;
    rd_mst_rdat_ready : out std_logic;
    rd_mst_rdat_data  : in  std_logic_vector(BUS_DATA_WIDTH-1 downto 0);
    rd_mst_rdat_last  : in  std_logic
  );
end entity;

architecture Implementation of Join_Mantle is
  component Join_Nucleus is
    generic (
      INDEX_WIDTH                    : integer := 32;
      TAG_WIDTH                      : integer := 1;
      SS_SOLD_DATE_SK_BUS_ADDR_WIDTH : integer := 64;
      SS_CDEMO_SK_BUS_ADDR_WIDTH     : integer := 64;
      SS_ADDR_SK_BUS_ADDR_WIDTH      : integer := 64;
      SS_STORE_SK_BUS_ADDR_WIDTH     : integer := 64;
      SS_QUANTITY_BUS_ADDR_WIDTH     : integer := 64;
      SS_SALES_PRICE_BUS_ADDR_WIDTH  : integer := 64;
      SS_NET_PROFIT_BUS_ADDR_WIDTH   : integer := 64
    );
    port (
      kcd_clk                      : in  std_logic;
      kcd_reset                    : in  std_logic;
      mmio_awvalid                 : in  std_logic;
      mmio_awready                 : out std_logic;
      mmio_awaddr                  : in  std_logic_vector(31 downto 0);
      mmio_wvalid                  : in  std_logic;
      mmio_wready                  : out std_logic;
      mmio_wdata                   : in  std_logic_vector(31 downto 0);
      mmio_wstrb                   : in  std_logic_vector(3 downto 0);
      mmio_bvalid                  : out std_logic;
      mmio_bready                  : in  std_logic;
      mmio_bresp                   : out std_logic_vector(1 downto 0);
      mmio_arvalid                 : in  std_logic;
      mmio_arready                 : out std_logic;
      mmio_araddr                  : in  std_logic_vector(31 downto 0);
      mmio_rvalid                  : out std_logic;
      mmio_rready                  : in  std_logic;
      mmio_rdata                   : out std_logic_vector(31 downto 0);
      mmio_rresp                   : out std_logic_vector(1 downto 0);
      ss_sold_date_sk_valid        : in  std_logic;
      ss_sold_date_sk_ready        : out std_logic;
      ss_sold_date_sk_dvalid       : in  std_logic;
      ss_sold_date_sk_last         : in  std_logic;
      ss_sold_date_sk              : in  std_logic_vector(63 downto 0);
      ss_cdemo_sk_valid            : in  std_logic;
      ss_cdemo_sk_ready            : out std_logic;
      ss_cdemo_sk_dvalid           : in  std_logic;
      ss_cdemo_sk_last             : in  std_logic;
      ss_cdemo_sk                  : in  std_logic_vector(63 downto 0);
      ss_addr_sk_valid             : in  std_logic;
      ss_addr_sk_ready             : out std_logic;
      ss_addr_sk_dvalid            : in  std_logic;
      ss_addr_sk_last              : in  std_logic;
      ss_addr_sk                   : in  std_logic_vector(63 downto 0);
      ss_store_sk_valid            : in  std_logic;
      ss_store_sk_ready            : out std_logic;
      ss_store_sk_dvalid           : in  std_logic;
      ss_store_sk_last             : in  std_logic;
      ss_store_sk                  : in  std_logic_vector(63 downto 0);
      ss_quantity_valid            : in  std_logic;
      ss_quantity_ready            : out std_logic;
      ss_quantity_dvalid           : in  std_logic;
      ss_quantity_last             : in  std_logic;
      ss_quantity                  : in  std_logic_vector(63 downto 0);
      ss_sales_price_valid         : in  std_logic;
      ss_sales_price_ready         : out std_logic;
      ss_sales_price_dvalid        : in  std_logic;
      ss_sales_price_last          : in  std_logic;
      ss_sales_price               : in  std_logic_vector(63 downto 0);
      ss_net_profit_valid          : in  std_logic;
      ss_net_profit_ready          : out std_logic;
      ss_net_profit_dvalid         : in  std_logic;
      ss_net_profit_last           : in  std_logic;
      ss_net_profit                : in  std_logic_vector(63 downto 0);
      ss_sold_date_sk_unl_valid    : in  std_logic;
      ss_sold_date_sk_unl_ready    : out std_logic;
      ss_sold_date_sk_unl_tag      : in  std_logic_vector(TAG_WIDTH-1 downto 0);
      ss_cdemo_sk_unl_valid        : in  std_logic;
      ss_cdemo_sk_unl_ready        : out std_logic;
      ss_cdemo_sk_unl_tag          : in  std_logic_vector(TAG_WIDTH-1 downto 0);
      ss_addr_sk_unl_valid         : in  std_logic;
      ss_addr_sk_unl_ready         : out std_logic;
      ss_addr_sk_unl_tag           : in  std_logic_vector(TAG_WIDTH-1 downto 0);
      ss_store_sk_unl_valid        : in  std_logic;
      ss_store_sk_unl_ready        : out std_logic;
      ss_store_sk_unl_tag          : in  std_logic_vector(TAG_WIDTH-1 downto 0);
      ss_quantity_unl_valid        : in  std_logic;
      ss_quantity_unl_ready        : out std_logic;
      ss_quantity_unl_tag          : in  std_logic_vector(TAG_WIDTH-1 downto 0);
      ss_sales_price_unl_valid     : in  std_logic;
      ss_sales_price_unl_ready     : out std_logic;
      ss_sales_price_unl_tag       : in  std_logic_vector(TAG_WIDTH-1 downto 0);
      ss_net_profit_unl_valid      : in  std_logic;
      ss_net_profit_unl_ready      : out std_logic;
      ss_net_profit_unl_tag        : in  std_logic_vector(TAG_WIDTH-1 downto 0);
      ss_sold_date_sk_cmd_valid    : out std_logic;
      ss_sold_date_sk_cmd_ready    : in  std_logic;
      ss_sold_date_sk_cmd_firstIdx : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      ss_sold_date_sk_cmd_lastIdx  : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      ss_sold_date_sk_cmd_ctrl     : out std_logic_vector(SS_SOLD_DATE_SK_BUS_ADDR_WIDTH-1 downto 0);
      ss_sold_date_sk_cmd_tag      : out std_logic_vector(TAG_WIDTH-1 downto 0);
      ss_cdemo_sk_cmd_valid        : out std_logic;
      ss_cdemo_sk_cmd_ready        : in  std_logic;
      ss_cdemo_sk_cmd_firstIdx     : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      ss_cdemo_sk_cmd_lastIdx      : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      ss_cdemo_sk_cmd_ctrl         : out std_logic_vector(SS_CDEMO_SK_BUS_ADDR_WIDTH-1 downto 0);
      ss_cdemo_sk_cmd_tag          : out std_logic_vector(TAG_WIDTH-1 downto 0);
      ss_addr_sk_cmd_valid         : out std_logic;
      ss_addr_sk_cmd_ready         : in  std_logic;
      ss_addr_sk_cmd_firstIdx      : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      ss_addr_sk_cmd_lastIdx       : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      ss_addr_sk_cmd_ctrl          : out std_logic_vector(SS_ADDR_SK_BUS_ADDR_WIDTH-1 downto 0);
      ss_addr_sk_cmd_tag           : out std_logic_vector(TAG_WIDTH-1 downto 0);
      ss_store_sk_cmd_valid        : out std_logic;
      ss_store_sk_cmd_ready        : in  std_logic;
      ss_store_sk_cmd_firstIdx     : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      ss_store_sk_cmd_lastIdx      : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      ss_store_sk_cmd_ctrl         : out std_logic_vector(SS_STORE_SK_BUS_ADDR_WIDTH-1 downto 0);
      ss_store_sk_cmd_tag          : out std_logic_vector(TAG_WIDTH-1 downto 0);
      ss_quantity_cmd_valid        : out std_logic;
      ss_quantity_cmd_ready        : in  std_logic;
      ss_quantity_cmd_firstIdx     : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      ss_quantity_cmd_lastIdx      : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      ss_quantity_cmd_ctrl         : out std_logic_vector(SS_QUANTITY_BUS_ADDR_WIDTH-1 downto 0);
      ss_quantity_cmd_tag          : out std_logic_vector(TAG_WIDTH-1 downto 0);
      ss_sales_price_cmd_valid     : out std_logic;
      ss_sales_price_cmd_ready     : in  std_logic;
      ss_sales_price_cmd_firstIdx  : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      ss_sales_price_cmd_lastIdx   : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      ss_sales_price_cmd_ctrl      : out std_logic_vector(SS_SALES_PRICE_BUS_ADDR_WIDTH-1 downto 0);
      ss_sales_price_cmd_tag       : out std_logic_vector(TAG_WIDTH-1 downto 0);
      ss_net_profit_cmd_valid      : out std_logic;
      ss_net_profit_cmd_ready      : in  std_logic;
      ss_net_profit_cmd_firstIdx   : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      ss_net_profit_cmd_lastIdx    : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      ss_net_profit_cmd_ctrl       : out std_logic_vector(SS_NET_PROFIT_BUS_ADDR_WIDTH-1 downto 0);
      ss_net_profit_cmd_tag        : out std_logic_vector(TAG_WIDTH-1 downto 0)
    );
  end component;

  component Join_ss is
    generic (
      INDEX_WIDTH                        : integer := 32;
      TAG_WIDTH                          : integer := 1;
      SS_SOLD_DATE_SK_BUS_ADDR_WIDTH     : integer := 64;
      SS_SOLD_DATE_SK_BUS_DATA_WIDTH     : integer := 512;
      SS_SOLD_DATE_SK_BUS_LEN_WIDTH      : integer := 8;
      SS_SOLD_DATE_SK_BUS_BURST_STEP_LEN : integer := 1;
      SS_SOLD_DATE_SK_BUS_BURST_MAX_LEN  : integer := 16;
      SS_CDEMO_SK_BUS_ADDR_WIDTH         : integer := 64;
      SS_CDEMO_SK_BUS_DATA_WIDTH         : integer := 512;
      SS_CDEMO_SK_BUS_LEN_WIDTH          : integer := 8;
      SS_CDEMO_SK_BUS_BURST_STEP_LEN     : integer := 1;
      SS_CDEMO_SK_BUS_BURST_MAX_LEN      : integer := 16;
      SS_ADDR_SK_BUS_ADDR_WIDTH          : integer := 64;
      SS_ADDR_SK_BUS_DATA_WIDTH          : integer := 512;
      SS_ADDR_SK_BUS_LEN_WIDTH           : integer := 8;
      SS_ADDR_SK_BUS_BURST_STEP_LEN      : integer := 1;
      SS_ADDR_SK_BUS_BURST_MAX_LEN       : integer := 16;
      SS_STORE_SK_BUS_ADDR_WIDTH         : integer := 64;
      SS_STORE_SK_BUS_DATA_WIDTH         : integer := 512;
      SS_STORE_SK_BUS_LEN_WIDTH          : integer := 8;
      SS_STORE_SK_BUS_BURST_STEP_LEN     : integer := 1;
      SS_STORE_SK_BUS_BURST_MAX_LEN      : integer := 16;
      SS_QUANTITY_BUS_ADDR_WIDTH         : integer := 64;
      SS_QUANTITY_BUS_DATA_WIDTH         : integer := 512;
      SS_QUANTITY_BUS_LEN_WIDTH          : integer := 8;
      SS_QUANTITY_BUS_BURST_STEP_LEN     : integer := 1;
      SS_QUANTITY_BUS_BURST_MAX_LEN      : integer := 16;
      SS_SALES_PRICE_BUS_ADDR_WIDTH      : integer := 64;
      SS_SALES_PRICE_BUS_DATA_WIDTH      : integer := 512;
      SS_SALES_PRICE_BUS_LEN_WIDTH       : integer := 8;
      SS_SALES_PRICE_BUS_BURST_STEP_LEN  : integer := 1;
      SS_SALES_PRICE_BUS_BURST_MAX_LEN   : integer := 16;
      SS_NET_PROFIT_BUS_ADDR_WIDTH       : integer := 64;
      SS_NET_PROFIT_BUS_DATA_WIDTH       : integer := 512;
      SS_NET_PROFIT_BUS_LEN_WIDTH        : integer := 8;
      SS_NET_PROFIT_BUS_BURST_STEP_LEN   : integer := 1;
      SS_NET_PROFIT_BUS_BURST_MAX_LEN    : integer := 16
    );
    port (
      bcd_clk                        : in  std_logic;
      bcd_reset                      : in  std_logic;
      kcd_clk                        : in  std_logic;
      kcd_reset                      : in  std_logic;
      ss_sold_date_sk_valid          : out std_logic;
      ss_sold_date_sk_ready          : in  std_logic;
      ss_sold_date_sk_dvalid         : out std_logic;
      ss_sold_date_sk_last           : out std_logic;
      ss_sold_date_sk                : out std_logic_vector(63 downto 0);
      ss_sold_date_sk_bus_rreq_valid : out std_logic;
      ss_sold_date_sk_bus_rreq_ready : in  std_logic;
      ss_sold_date_sk_bus_rreq_addr  : out std_logic_vector(SS_SOLD_DATE_SK_BUS_ADDR_WIDTH-1 downto 0);
      ss_sold_date_sk_bus_rreq_len   : out std_logic_vector(SS_SOLD_DATE_SK_BUS_LEN_WIDTH-1 downto 0);
      ss_sold_date_sk_bus_rdat_valid : in  std_logic;
      ss_sold_date_sk_bus_rdat_ready : out std_logic;
      ss_sold_date_sk_bus_rdat_data  : in  std_logic_vector(SS_SOLD_DATE_SK_BUS_DATA_WIDTH-1 downto 0);
      ss_sold_date_sk_bus_rdat_last  : in  std_logic;
      ss_sold_date_sk_cmd_valid      : in  std_logic;
      ss_sold_date_sk_cmd_ready      : out std_logic;
      ss_sold_date_sk_cmd_firstIdx   : in  std_logic_vector(INDEX_WIDTH-1 downto 0);
      ss_sold_date_sk_cmd_lastIdx    : in  std_logic_vector(INDEX_WIDTH-1 downto 0);
      ss_sold_date_sk_cmd_ctrl       : in  std_logic_vector(SS_SOLD_DATE_SK_BUS_ADDR_WIDTH-1 downto 0);
      ss_sold_date_sk_cmd_tag        : in  std_logic_vector(TAG_WIDTH-1 downto 0);
      ss_sold_date_sk_unl_valid      : out std_logic;
      ss_sold_date_sk_unl_ready      : in  std_logic;
      ss_sold_date_sk_unl_tag        : out std_logic_vector(TAG_WIDTH-1 downto 0);
      ss_cdemo_sk_valid              : out std_logic;
      ss_cdemo_sk_ready              : in  std_logic;
      ss_cdemo_sk_dvalid             : out std_logic;
      ss_cdemo_sk_last               : out std_logic;
      ss_cdemo_sk                    : out std_logic_vector(63 downto 0);
      ss_cdemo_sk_bus_rreq_valid     : out std_logic;
      ss_cdemo_sk_bus_rreq_ready     : in  std_logic;
      ss_cdemo_sk_bus_rreq_addr      : out std_logic_vector(SS_CDEMO_SK_BUS_ADDR_WIDTH-1 downto 0);
      ss_cdemo_sk_bus_rreq_len       : out std_logic_vector(SS_CDEMO_SK_BUS_LEN_WIDTH-1 downto 0);
      ss_cdemo_sk_bus_rdat_valid     : in  std_logic;
      ss_cdemo_sk_bus_rdat_ready     : out std_logic;
      ss_cdemo_sk_bus_rdat_data      : in  std_logic_vector(SS_CDEMO_SK_BUS_DATA_WIDTH-1 downto 0);
      ss_cdemo_sk_bus_rdat_last      : in  std_logic;
      ss_cdemo_sk_cmd_valid          : in  std_logic;
      ss_cdemo_sk_cmd_ready          : out std_logic;
      ss_cdemo_sk_cmd_firstIdx       : in  std_logic_vector(INDEX_WIDTH-1 downto 0);
      ss_cdemo_sk_cmd_lastIdx        : in  std_logic_vector(INDEX_WIDTH-1 downto 0);
      ss_cdemo_sk_cmd_ctrl           : in  std_logic_vector(SS_CDEMO_SK_BUS_ADDR_WIDTH-1 downto 0);
      ss_cdemo_sk_cmd_tag            : in  std_logic_vector(TAG_WIDTH-1 downto 0);
      ss_cdemo_sk_unl_valid          : out std_logic;
      ss_cdemo_sk_unl_ready          : in  std_logic;
      ss_cdemo_sk_unl_tag            : out std_logic_vector(TAG_WIDTH-1 downto 0);
      ss_addr_sk_valid               : out std_logic;
      ss_addr_sk_ready               : in  std_logic;
      ss_addr_sk_dvalid              : out std_logic;
      ss_addr_sk_last                : out std_logic;
      ss_addr_sk                     : out std_logic_vector(63 downto 0);
      ss_addr_sk_bus_rreq_valid      : out std_logic;
      ss_addr_sk_bus_rreq_ready      : in  std_logic;
      ss_addr_sk_bus_rreq_addr       : out std_logic_vector(SS_ADDR_SK_BUS_ADDR_WIDTH-1 downto 0);
      ss_addr_sk_bus_rreq_len        : out std_logic_vector(SS_ADDR_SK_BUS_LEN_WIDTH-1 downto 0);
      ss_addr_sk_bus_rdat_valid      : in  std_logic;
      ss_addr_sk_bus_rdat_ready      : out std_logic;
      ss_addr_sk_bus_rdat_data       : in  std_logic_vector(SS_ADDR_SK_BUS_DATA_WIDTH-1 downto 0);
      ss_addr_sk_bus_rdat_last       : in  std_logic;
      ss_addr_sk_cmd_valid           : in  std_logic;
      ss_addr_sk_cmd_ready           : out std_logic;
      ss_addr_sk_cmd_firstIdx        : in  std_logic_vector(INDEX_WIDTH-1 downto 0);
      ss_addr_sk_cmd_lastIdx         : in  std_logic_vector(INDEX_WIDTH-1 downto 0);
      ss_addr_sk_cmd_ctrl            : in  std_logic_vector(SS_ADDR_SK_BUS_ADDR_WIDTH-1 downto 0);
      ss_addr_sk_cmd_tag             : in  std_logic_vector(TAG_WIDTH-1 downto 0);
      ss_addr_sk_unl_valid           : out std_logic;
      ss_addr_sk_unl_ready           : in  std_logic;
      ss_addr_sk_unl_tag             : out std_logic_vector(TAG_WIDTH-1 downto 0);
      ss_store_sk_valid              : out std_logic;
      ss_store_sk_ready              : in  std_logic;
      ss_store_sk_dvalid             : out std_logic;
      ss_store_sk_last               : out std_logic;
      ss_store_sk                    : out std_logic_vector(63 downto 0);
      ss_store_sk_bus_rreq_valid     : out std_logic;
      ss_store_sk_bus_rreq_ready     : in  std_logic;
      ss_store_sk_bus_rreq_addr      : out std_logic_vector(SS_STORE_SK_BUS_ADDR_WIDTH-1 downto 0);
      ss_store_sk_bus_rreq_len       : out std_logic_vector(SS_STORE_SK_BUS_LEN_WIDTH-1 downto 0);
      ss_store_sk_bus_rdat_valid     : in  std_logic;
      ss_store_sk_bus_rdat_ready     : out std_logic;
      ss_store_sk_bus_rdat_data      : in  std_logic_vector(SS_STORE_SK_BUS_DATA_WIDTH-1 downto 0);
      ss_store_sk_bus_rdat_last      : in  std_logic;
      ss_store_sk_cmd_valid          : in  std_logic;
      ss_store_sk_cmd_ready          : out std_logic;
      ss_store_sk_cmd_firstIdx       : in  std_logic_vector(INDEX_WIDTH-1 downto 0);
      ss_store_sk_cmd_lastIdx        : in  std_logic_vector(INDEX_WIDTH-1 downto 0);
      ss_store_sk_cmd_ctrl           : in  std_logic_vector(SS_STORE_SK_BUS_ADDR_WIDTH-1 downto 0);
      ss_store_sk_cmd_tag            : in  std_logic_vector(TAG_WIDTH-1 downto 0);
      ss_store_sk_unl_valid          : out std_logic;
      ss_store_sk_unl_ready          : in  std_logic;
      ss_store_sk_unl_tag            : out std_logic_vector(TAG_WIDTH-1 downto 0);
      ss_quantity_valid              : out std_logic;
      ss_quantity_ready              : in  std_logic;
      ss_quantity_dvalid             : out std_logic;
      ss_quantity_last               : out std_logic;
      ss_quantity                    : out std_logic_vector(63 downto 0);
      ss_quantity_bus_rreq_valid     : out std_logic;
      ss_quantity_bus_rreq_ready     : in  std_logic;
      ss_quantity_bus_rreq_addr      : out std_logic_vector(SS_QUANTITY_BUS_ADDR_WIDTH-1 downto 0);
      ss_quantity_bus_rreq_len       : out std_logic_vector(SS_QUANTITY_BUS_LEN_WIDTH-1 downto 0);
      ss_quantity_bus_rdat_valid     : in  std_logic;
      ss_quantity_bus_rdat_ready     : out std_logic;
      ss_quantity_bus_rdat_data      : in  std_logic_vector(SS_QUANTITY_BUS_DATA_WIDTH-1 downto 0);
      ss_quantity_bus_rdat_last      : in  std_logic;
      ss_quantity_cmd_valid          : in  std_logic;
      ss_quantity_cmd_ready          : out std_logic;
      ss_quantity_cmd_firstIdx       : in  std_logic_vector(INDEX_WIDTH-1 downto 0);
      ss_quantity_cmd_lastIdx        : in  std_logic_vector(INDEX_WIDTH-1 downto 0);
      ss_quantity_cmd_ctrl           : in  std_logic_vector(SS_QUANTITY_BUS_ADDR_WIDTH-1 downto 0);
      ss_quantity_cmd_tag            : in  std_logic_vector(TAG_WIDTH-1 downto 0);
      ss_quantity_unl_valid          : out std_logic;
      ss_quantity_unl_ready          : in  std_logic;
      ss_quantity_unl_tag            : out std_logic_vector(TAG_WIDTH-1 downto 0);
      ss_sales_price_valid           : out std_logic;
      ss_sales_price_ready           : in  std_logic;
      ss_sales_price_dvalid          : out std_logic;
      ss_sales_price_last            : out std_logic;
      ss_sales_price                 : out std_logic_vector(63 downto 0);
      ss_sales_price_bus_rreq_valid  : out std_logic;
      ss_sales_price_bus_rreq_ready  : in  std_logic;
      ss_sales_price_bus_rreq_addr   : out std_logic_vector(SS_SALES_PRICE_BUS_ADDR_WIDTH-1 downto 0);
      ss_sales_price_bus_rreq_len    : out std_logic_vector(SS_SALES_PRICE_BUS_LEN_WIDTH-1 downto 0);
      ss_sales_price_bus_rdat_valid  : in  std_logic;
      ss_sales_price_bus_rdat_ready  : out std_logic;
      ss_sales_price_bus_rdat_data   : in  std_logic_vector(SS_SALES_PRICE_BUS_DATA_WIDTH-1 downto 0);
      ss_sales_price_bus_rdat_last   : in  std_logic;
      ss_sales_price_cmd_valid       : in  std_logic;
      ss_sales_price_cmd_ready       : out std_logic;
      ss_sales_price_cmd_firstIdx    : in  std_logic_vector(INDEX_WIDTH-1 downto 0);
      ss_sales_price_cmd_lastIdx     : in  std_logic_vector(INDEX_WIDTH-1 downto 0);
      ss_sales_price_cmd_ctrl        : in  std_logic_vector(SS_SALES_PRICE_BUS_ADDR_WIDTH-1 downto 0);
      ss_sales_price_cmd_tag         : in  std_logic_vector(TAG_WIDTH-1 downto 0);
      ss_sales_price_unl_valid       : out std_logic;
      ss_sales_price_unl_ready       : in  std_logic;
      ss_sales_price_unl_tag         : out std_logic_vector(TAG_WIDTH-1 downto 0);
      ss_net_profit_valid            : out std_logic;
      ss_net_profit_ready            : in  std_logic;
      ss_net_profit_dvalid           : out std_logic;
      ss_net_profit_last             : out std_logic;
      ss_net_profit                  : out std_logic_vector(63 downto 0);
      ss_net_profit_bus_rreq_valid   : out std_logic;
      ss_net_profit_bus_rreq_ready   : in  std_logic;
      ss_net_profit_bus_rreq_addr    : out std_logic_vector(SS_NET_PROFIT_BUS_ADDR_WIDTH-1 downto 0);
      ss_net_profit_bus_rreq_len     : out std_logic_vector(SS_NET_PROFIT_BUS_LEN_WIDTH-1 downto 0);
      ss_net_profit_bus_rdat_valid   : in  std_logic;
      ss_net_profit_bus_rdat_ready   : out std_logic;
      ss_net_profit_bus_rdat_data    : in  std_logic_vector(SS_NET_PROFIT_BUS_DATA_WIDTH-1 downto 0);
      ss_net_profit_bus_rdat_last    : in  std_logic;
      ss_net_profit_cmd_valid        : in  std_logic;
      ss_net_profit_cmd_ready        : out std_logic;
      ss_net_profit_cmd_firstIdx     : in  std_logic_vector(INDEX_WIDTH-1 downto 0);
      ss_net_profit_cmd_lastIdx      : in  std_logic_vector(INDEX_WIDTH-1 downto 0);
      ss_net_profit_cmd_ctrl         : in  std_logic_vector(SS_NET_PROFIT_BUS_ADDR_WIDTH-1 downto 0);
      ss_net_profit_cmd_tag          : in  std_logic_vector(TAG_WIDTH-1 downto 0);
      ss_net_profit_unl_valid        : out std_logic;
      ss_net_profit_unl_ready        : in  std_logic;
      ss_net_profit_unl_tag          : out std_logic_vector(TAG_WIDTH-1 downto 0)
    );
  end component;

  signal Join_Nucleus_inst_mmio_awvalid                 : std_logic;
  signal Join_Nucleus_inst_mmio_awready                 : std_logic;
  signal Join_Nucleus_inst_mmio_awaddr                  : std_logic_vector(31 downto 0);
  signal Join_Nucleus_inst_mmio_wvalid                  : std_logic;
  signal Join_Nucleus_inst_mmio_wready                  : std_logic;
  signal Join_Nucleus_inst_mmio_wdata                   : std_logic_vector(31 downto 0);
  signal Join_Nucleus_inst_mmio_wstrb                   : std_logic_vector(3 downto 0);
  signal Join_Nucleus_inst_mmio_bvalid                  : std_logic;
  signal Join_Nucleus_inst_mmio_bready                  : std_logic;
  signal Join_Nucleus_inst_mmio_bresp                   : std_logic_vector(1 downto 0);
  signal Join_Nucleus_inst_mmio_arvalid                 : std_logic;
  signal Join_Nucleus_inst_mmio_arready                 : std_logic;
  signal Join_Nucleus_inst_mmio_araddr                  : std_logic_vector(31 downto 0);
  signal Join_Nucleus_inst_mmio_rvalid                  : std_logic;
  signal Join_Nucleus_inst_mmio_rready                  : std_logic;
  signal Join_Nucleus_inst_mmio_rdata                   : std_logic_vector(31 downto 0);
  signal Join_Nucleus_inst_mmio_rresp                   : std_logic_vector(1 downto 0);

  signal Join_Nucleus_inst_ss_sold_date_sk_valid        : std_logic;
  signal Join_Nucleus_inst_ss_sold_date_sk_ready        : std_logic;
  signal Join_Nucleus_inst_ss_sold_date_sk_dvalid       : std_logic;
  signal Join_Nucleus_inst_ss_sold_date_sk_last         : std_logic;
  signal Join_Nucleus_inst_ss_sold_date_sk              : std_logic_vector(63 downto 0);

  signal Join_Nucleus_inst_ss_cdemo_sk_valid            : std_logic;
  signal Join_Nucleus_inst_ss_cdemo_sk_ready            : std_logic;
  signal Join_Nucleus_inst_ss_cdemo_sk_dvalid           : std_logic;
  signal Join_Nucleus_inst_ss_cdemo_sk_last             : std_logic;
  signal Join_Nucleus_inst_ss_cdemo_sk                  : std_logic_vector(63 downto 0);

  signal Join_Nucleus_inst_ss_addr_sk_valid             : std_logic;
  signal Join_Nucleus_inst_ss_addr_sk_ready             : std_logic;
  signal Join_Nucleus_inst_ss_addr_sk_dvalid            : std_logic;
  signal Join_Nucleus_inst_ss_addr_sk_last              : std_logic;
  signal Join_Nucleus_inst_ss_addr_sk                   : std_logic_vector(63 downto 0);

  signal Join_Nucleus_inst_ss_store_sk_valid            : std_logic;
  signal Join_Nucleus_inst_ss_store_sk_ready            : std_logic;
  signal Join_Nucleus_inst_ss_store_sk_dvalid           : std_logic;
  signal Join_Nucleus_inst_ss_store_sk_last             : std_logic;
  signal Join_Nucleus_inst_ss_store_sk                  : std_logic_vector(63 downto 0);

  signal Join_Nucleus_inst_ss_quantity_valid            : std_logic;
  signal Join_Nucleus_inst_ss_quantity_ready            : std_logic;
  signal Join_Nucleus_inst_ss_quantity_dvalid           : std_logic;
  signal Join_Nucleus_inst_ss_quantity_last             : std_logic;
  signal Join_Nucleus_inst_ss_quantity                  : std_logic_vector(63 downto 0);

  signal Join_Nucleus_inst_ss_sales_price_valid         : std_logic;
  signal Join_Nucleus_inst_ss_sales_price_ready         : std_logic;
  signal Join_Nucleus_inst_ss_sales_price_dvalid        : std_logic;
  signal Join_Nucleus_inst_ss_sales_price_last          : std_logic;
  signal Join_Nucleus_inst_ss_sales_price               : std_logic_vector(63 downto 0);

  signal Join_Nucleus_inst_ss_net_profit_valid          : std_logic;
  signal Join_Nucleus_inst_ss_net_profit_ready          : std_logic;
  signal Join_Nucleus_inst_ss_net_profit_dvalid         : std_logic;
  signal Join_Nucleus_inst_ss_net_profit_last           : std_logic;
  signal Join_Nucleus_inst_ss_net_profit                : std_logic_vector(63 downto 0);

  signal Join_Nucleus_inst_ss_sold_date_sk_unl_valid    : std_logic;
  signal Join_Nucleus_inst_ss_sold_date_sk_unl_ready    : std_logic;
  signal Join_Nucleus_inst_ss_sold_date_sk_unl_tag      : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal Join_Nucleus_inst_ss_cdemo_sk_unl_valid        : std_logic;
  signal Join_Nucleus_inst_ss_cdemo_sk_unl_ready        : std_logic;
  signal Join_Nucleus_inst_ss_cdemo_sk_unl_tag          : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal Join_Nucleus_inst_ss_addr_sk_unl_valid         : std_logic;
  signal Join_Nucleus_inst_ss_addr_sk_unl_ready         : std_logic;
  signal Join_Nucleus_inst_ss_addr_sk_unl_tag           : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal Join_Nucleus_inst_ss_store_sk_unl_valid        : std_logic;
  signal Join_Nucleus_inst_ss_store_sk_unl_ready        : std_logic;
  signal Join_Nucleus_inst_ss_store_sk_unl_tag          : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal Join_Nucleus_inst_ss_quantity_unl_valid        : std_logic;
  signal Join_Nucleus_inst_ss_quantity_unl_ready        : std_logic;
  signal Join_Nucleus_inst_ss_quantity_unl_tag          : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal Join_Nucleus_inst_ss_sales_price_unl_valid     : std_logic;
  signal Join_Nucleus_inst_ss_sales_price_unl_ready     : std_logic;
  signal Join_Nucleus_inst_ss_sales_price_unl_tag       : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal Join_Nucleus_inst_ss_net_profit_unl_valid      : std_logic;
  signal Join_Nucleus_inst_ss_net_profit_unl_ready      : std_logic;
  signal Join_Nucleus_inst_ss_net_profit_unl_tag        : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal Join_Nucleus_inst_ss_sold_date_sk_cmd_valid    : std_logic;
  signal Join_Nucleus_inst_ss_sold_date_sk_cmd_ready    : std_logic;
  signal Join_Nucleus_inst_ss_sold_date_sk_cmd_firstIdx : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal Join_Nucleus_inst_ss_sold_date_sk_cmd_lastIdx  : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal Join_Nucleus_inst_ss_sold_date_sk_cmd_ctrl     : std_logic_vector(BUS_ADDR_WIDTH-1 downto 0);
  signal Join_Nucleus_inst_ss_sold_date_sk_cmd_tag      : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal Join_Nucleus_inst_ss_cdemo_sk_cmd_valid        : std_logic;
  signal Join_Nucleus_inst_ss_cdemo_sk_cmd_ready        : std_logic;
  signal Join_Nucleus_inst_ss_cdemo_sk_cmd_firstIdx     : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal Join_Nucleus_inst_ss_cdemo_sk_cmd_lastIdx      : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal Join_Nucleus_inst_ss_cdemo_sk_cmd_ctrl         : std_logic_vector(BUS_ADDR_WIDTH-1 downto 0);
  signal Join_Nucleus_inst_ss_cdemo_sk_cmd_tag          : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal Join_Nucleus_inst_ss_addr_sk_cmd_valid         : std_logic;
  signal Join_Nucleus_inst_ss_addr_sk_cmd_ready         : std_logic;
  signal Join_Nucleus_inst_ss_addr_sk_cmd_firstIdx      : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal Join_Nucleus_inst_ss_addr_sk_cmd_lastIdx       : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal Join_Nucleus_inst_ss_addr_sk_cmd_ctrl          : std_logic_vector(BUS_ADDR_WIDTH-1 downto 0);
  signal Join_Nucleus_inst_ss_addr_sk_cmd_tag           : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal Join_Nucleus_inst_ss_store_sk_cmd_valid        : std_logic;
  signal Join_Nucleus_inst_ss_store_sk_cmd_ready        : std_logic;
  signal Join_Nucleus_inst_ss_store_sk_cmd_firstIdx     : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal Join_Nucleus_inst_ss_store_sk_cmd_lastIdx      : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal Join_Nucleus_inst_ss_store_sk_cmd_ctrl         : std_logic_vector(BUS_ADDR_WIDTH-1 downto 0);
  signal Join_Nucleus_inst_ss_store_sk_cmd_tag          : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal Join_Nucleus_inst_ss_quantity_cmd_valid        : std_logic;
  signal Join_Nucleus_inst_ss_quantity_cmd_ready        : std_logic;
  signal Join_Nucleus_inst_ss_quantity_cmd_firstIdx     : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal Join_Nucleus_inst_ss_quantity_cmd_lastIdx      : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal Join_Nucleus_inst_ss_quantity_cmd_ctrl         : std_logic_vector(BUS_ADDR_WIDTH-1 downto 0);
  signal Join_Nucleus_inst_ss_quantity_cmd_tag          : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal Join_Nucleus_inst_ss_sales_price_cmd_valid     : std_logic;
  signal Join_Nucleus_inst_ss_sales_price_cmd_ready     : std_logic;
  signal Join_Nucleus_inst_ss_sales_price_cmd_firstIdx  : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal Join_Nucleus_inst_ss_sales_price_cmd_lastIdx   : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal Join_Nucleus_inst_ss_sales_price_cmd_ctrl      : std_logic_vector(BUS_ADDR_WIDTH-1 downto 0);
  signal Join_Nucleus_inst_ss_sales_price_cmd_tag       : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal Join_Nucleus_inst_ss_net_profit_cmd_valid      : std_logic;
  signal Join_Nucleus_inst_ss_net_profit_cmd_ready      : std_logic;
  signal Join_Nucleus_inst_ss_net_profit_cmd_firstIdx   : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal Join_Nucleus_inst_ss_net_profit_cmd_lastIdx    : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal Join_Nucleus_inst_ss_net_profit_cmd_ctrl       : std_logic_vector(BUS_ADDR_WIDTH-1 downto 0);
  signal Join_Nucleus_inst_ss_net_profit_cmd_tag        : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal Join_ss_inst_ss_sold_date_sk_valid             : std_logic;
  signal Join_ss_inst_ss_sold_date_sk_ready             : std_logic;
  signal Join_ss_inst_ss_sold_date_sk_dvalid            : std_logic;
  signal Join_ss_inst_ss_sold_date_sk_last              : std_logic;
  signal Join_ss_inst_ss_sold_date_sk                   : std_logic_vector(63 downto 0);

  signal Join_ss_inst_ss_sold_date_sk_bus_rreq_valid    : std_logic;
  signal Join_ss_inst_ss_sold_date_sk_bus_rreq_ready    : std_logic;
  signal Join_ss_inst_ss_sold_date_sk_bus_rreq_addr     : std_logic_vector(BUS_ADDR_WIDTH-1 downto 0);
  signal Join_ss_inst_ss_sold_date_sk_bus_rreq_len      : std_logic_vector(BUS_LEN_WIDTH-1 downto 0);
  signal Join_ss_inst_ss_sold_date_sk_bus_rdat_valid    : std_logic;
  signal Join_ss_inst_ss_sold_date_sk_bus_rdat_ready    : std_logic;
  signal Join_ss_inst_ss_sold_date_sk_bus_rdat_data     : std_logic_vector(BUS_DATA_WIDTH-1 downto 0);
  signal Join_ss_inst_ss_sold_date_sk_bus_rdat_last     : std_logic;

  signal Join_ss_inst_ss_sold_date_sk_cmd_valid         : std_logic;
  signal Join_ss_inst_ss_sold_date_sk_cmd_ready         : std_logic;
  signal Join_ss_inst_ss_sold_date_sk_cmd_firstIdx      : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal Join_ss_inst_ss_sold_date_sk_cmd_lastIdx       : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal Join_ss_inst_ss_sold_date_sk_cmd_ctrl          : std_logic_vector(BUS_ADDR_WIDTH-1 downto 0);
  signal Join_ss_inst_ss_sold_date_sk_cmd_tag           : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal Join_ss_inst_ss_sold_date_sk_unl_valid         : std_logic;
  signal Join_ss_inst_ss_sold_date_sk_unl_ready         : std_logic;
  signal Join_ss_inst_ss_sold_date_sk_unl_tag           : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal Join_ss_inst_ss_cdemo_sk_valid                 : std_logic;
  signal Join_ss_inst_ss_cdemo_sk_ready                 : std_logic;
  signal Join_ss_inst_ss_cdemo_sk_dvalid                : std_logic;
  signal Join_ss_inst_ss_cdemo_sk_last                  : std_logic;
  signal Join_ss_inst_ss_cdemo_sk                       : std_logic_vector(63 downto 0);

  signal Join_ss_inst_ss_cdemo_sk_bus_rreq_valid        : std_logic;
  signal Join_ss_inst_ss_cdemo_sk_bus_rreq_ready        : std_logic;
  signal Join_ss_inst_ss_cdemo_sk_bus_rreq_addr         : std_logic_vector(BUS_ADDR_WIDTH-1 downto 0);
  signal Join_ss_inst_ss_cdemo_sk_bus_rreq_len          : std_logic_vector(BUS_LEN_WIDTH-1 downto 0);
  signal Join_ss_inst_ss_cdemo_sk_bus_rdat_valid        : std_logic;
  signal Join_ss_inst_ss_cdemo_sk_bus_rdat_ready        : std_logic;
  signal Join_ss_inst_ss_cdemo_sk_bus_rdat_data         : std_logic_vector(BUS_DATA_WIDTH-1 downto 0);
  signal Join_ss_inst_ss_cdemo_sk_bus_rdat_last         : std_logic;

  signal Join_ss_inst_ss_cdemo_sk_cmd_valid             : std_logic;
  signal Join_ss_inst_ss_cdemo_sk_cmd_ready             : std_logic;
  signal Join_ss_inst_ss_cdemo_sk_cmd_firstIdx          : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal Join_ss_inst_ss_cdemo_sk_cmd_lastIdx           : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal Join_ss_inst_ss_cdemo_sk_cmd_ctrl              : std_logic_vector(BUS_ADDR_WIDTH-1 downto 0);
  signal Join_ss_inst_ss_cdemo_sk_cmd_tag               : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal Join_ss_inst_ss_cdemo_sk_unl_valid             : std_logic;
  signal Join_ss_inst_ss_cdemo_sk_unl_ready             : std_logic;
  signal Join_ss_inst_ss_cdemo_sk_unl_tag               : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal Join_ss_inst_ss_addr_sk_valid                  : std_logic;
  signal Join_ss_inst_ss_addr_sk_ready                  : std_logic;
  signal Join_ss_inst_ss_addr_sk_dvalid                 : std_logic;
  signal Join_ss_inst_ss_addr_sk_last                   : std_logic;
  signal Join_ss_inst_ss_addr_sk                        : std_logic_vector(63 downto 0);

  signal Join_ss_inst_ss_addr_sk_bus_rreq_valid         : std_logic;
  signal Join_ss_inst_ss_addr_sk_bus_rreq_ready         : std_logic;
  signal Join_ss_inst_ss_addr_sk_bus_rreq_addr          : std_logic_vector(BUS_ADDR_WIDTH-1 downto 0);
  signal Join_ss_inst_ss_addr_sk_bus_rreq_len           : std_logic_vector(BUS_LEN_WIDTH-1 downto 0);
  signal Join_ss_inst_ss_addr_sk_bus_rdat_valid         : std_logic;
  signal Join_ss_inst_ss_addr_sk_bus_rdat_ready         : std_logic;
  signal Join_ss_inst_ss_addr_sk_bus_rdat_data          : std_logic_vector(BUS_DATA_WIDTH-1 downto 0);
  signal Join_ss_inst_ss_addr_sk_bus_rdat_last          : std_logic;

  signal Join_ss_inst_ss_addr_sk_cmd_valid              : std_logic;
  signal Join_ss_inst_ss_addr_sk_cmd_ready              : std_logic;
  signal Join_ss_inst_ss_addr_sk_cmd_firstIdx           : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal Join_ss_inst_ss_addr_sk_cmd_lastIdx            : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal Join_ss_inst_ss_addr_sk_cmd_ctrl               : std_logic_vector(BUS_ADDR_WIDTH-1 downto 0);
  signal Join_ss_inst_ss_addr_sk_cmd_tag                : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal Join_ss_inst_ss_addr_sk_unl_valid              : std_logic;
  signal Join_ss_inst_ss_addr_sk_unl_ready              : std_logic;
  signal Join_ss_inst_ss_addr_sk_unl_tag                : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal Join_ss_inst_ss_store_sk_valid                 : std_logic;
  signal Join_ss_inst_ss_store_sk_ready                 : std_logic;
  signal Join_ss_inst_ss_store_sk_dvalid                : std_logic;
  signal Join_ss_inst_ss_store_sk_last                  : std_logic;
  signal Join_ss_inst_ss_store_sk                       : std_logic_vector(63 downto 0);

  signal Join_ss_inst_ss_store_sk_bus_rreq_valid        : std_logic;
  signal Join_ss_inst_ss_store_sk_bus_rreq_ready        : std_logic;
  signal Join_ss_inst_ss_store_sk_bus_rreq_addr         : std_logic_vector(BUS_ADDR_WIDTH-1 downto 0);
  signal Join_ss_inst_ss_store_sk_bus_rreq_len          : std_logic_vector(BUS_LEN_WIDTH-1 downto 0);
  signal Join_ss_inst_ss_store_sk_bus_rdat_valid        : std_logic;
  signal Join_ss_inst_ss_store_sk_bus_rdat_ready        : std_logic;
  signal Join_ss_inst_ss_store_sk_bus_rdat_data         : std_logic_vector(BUS_DATA_WIDTH-1 downto 0);
  signal Join_ss_inst_ss_store_sk_bus_rdat_last         : std_logic;

  signal Join_ss_inst_ss_store_sk_cmd_valid             : std_logic;
  signal Join_ss_inst_ss_store_sk_cmd_ready             : std_logic;
  signal Join_ss_inst_ss_store_sk_cmd_firstIdx          : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal Join_ss_inst_ss_store_sk_cmd_lastIdx           : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal Join_ss_inst_ss_store_sk_cmd_ctrl              : std_logic_vector(BUS_ADDR_WIDTH-1 downto 0);
  signal Join_ss_inst_ss_store_sk_cmd_tag               : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal Join_ss_inst_ss_store_sk_unl_valid             : std_logic;
  signal Join_ss_inst_ss_store_sk_unl_ready             : std_logic;
  signal Join_ss_inst_ss_store_sk_unl_tag               : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal Join_ss_inst_ss_quantity_valid                 : std_logic;
  signal Join_ss_inst_ss_quantity_ready                 : std_logic;
  signal Join_ss_inst_ss_quantity_dvalid                : std_logic;
  signal Join_ss_inst_ss_quantity_last                  : std_logic;
  signal Join_ss_inst_ss_quantity                       : std_logic_vector(63 downto 0);

  signal Join_ss_inst_ss_quantity_bus_rreq_valid        : std_logic;
  signal Join_ss_inst_ss_quantity_bus_rreq_ready        : std_logic;
  signal Join_ss_inst_ss_quantity_bus_rreq_addr         : std_logic_vector(BUS_ADDR_WIDTH-1 downto 0);
  signal Join_ss_inst_ss_quantity_bus_rreq_len          : std_logic_vector(BUS_LEN_WIDTH-1 downto 0);
  signal Join_ss_inst_ss_quantity_bus_rdat_valid        : std_logic;
  signal Join_ss_inst_ss_quantity_bus_rdat_ready        : std_logic;
  signal Join_ss_inst_ss_quantity_bus_rdat_data         : std_logic_vector(BUS_DATA_WIDTH-1 downto 0);
  signal Join_ss_inst_ss_quantity_bus_rdat_last         : std_logic;

  signal Join_ss_inst_ss_quantity_cmd_valid             : std_logic;
  signal Join_ss_inst_ss_quantity_cmd_ready             : std_logic;
  signal Join_ss_inst_ss_quantity_cmd_firstIdx          : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal Join_ss_inst_ss_quantity_cmd_lastIdx           : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal Join_ss_inst_ss_quantity_cmd_ctrl              : std_logic_vector(BUS_ADDR_WIDTH-1 downto 0);
  signal Join_ss_inst_ss_quantity_cmd_tag               : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal Join_ss_inst_ss_quantity_unl_valid             : std_logic;
  signal Join_ss_inst_ss_quantity_unl_ready             : std_logic;
  signal Join_ss_inst_ss_quantity_unl_tag               : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal Join_ss_inst_ss_sales_price_valid              : std_logic;
  signal Join_ss_inst_ss_sales_price_ready              : std_logic;
  signal Join_ss_inst_ss_sales_price_dvalid             : std_logic;
  signal Join_ss_inst_ss_sales_price_last               : std_logic;
  signal Join_ss_inst_ss_sales_price                    : std_logic_vector(63 downto 0);

  signal Join_ss_inst_ss_sales_price_bus_rreq_valid     : std_logic;
  signal Join_ss_inst_ss_sales_price_bus_rreq_ready     : std_logic;
  signal Join_ss_inst_ss_sales_price_bus_rreq_addr      : std_logic_vector(BUS_ADDR_WIDTH-1 downto 0);
  signal Join_ss_inst_ss_sales_price_bus_rreq_len       : std_logic_vector(BUS_LEN_WIDTH-1 downto 0);
  signal Join_ss_inst_ss_sales_price_bus_rdat_valid     : std_logic;
  signal Join_ss_inst_ss_sales_price_bus_rdat_ready     : std_logic;
  signal Join_ss_inst_ss_sales_price_bus_rdat_data      : std_logic_vector(BUS_DATA_WIDTH-1 downto 0);
  signal Join_ss_inst_ss_sales_price_bus_rdat_last      : std_logic;

  signal Join_ss_inst_ss_sales_price_cmd_valid          : std_logic;
  signal Join_ss_inst_ss_sales_price_cmd_ready          : std_logic;
  signal Join_ss_inst_ss_sales_price_cmd_firstIdx       : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal Join_ss_inst_ss_sales_price_cmd_lastIdx        : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal Join_ss_inst_ss_sales_price_cmd_ctrl           : std_logic_vector(BUS_ADDR_WIDTH-1 downto 0);
  signal Join_ss_inst_ss_sales_price_cmd_tag            : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal Join_ss_inst_ss_sales_price_unl_valid          : std_logic;
  signal Join_ss_inst_ss_sales_price_unl_ready          : std_logic;
  signal Join_ss_inst_ss_sales_price_unl_tag            : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal Join_ss_inst_ss_net_profit_valid               : std_logic;
  signal Join_ss_inst_ss_net_profit_ready               : std_logic;
  signal Join_ss_inst_ss_net_profit_dvalid              : std_logic;
  signal Join_ss_inst_ss_net_profit_last                : std_logic;
  signal Join_ss_inst_ss_net_profit                     : std_logic_vector(63 downto 0);

  signal Join_ss_inst_ss_net_profit_bus_rreq_valid      : std_logic;
  signal Join_ss_inst_ss_net_profit_bus_rreq_ready      : std_logic;
  signal Join_ss_inst_ss_net_profit_bus_rreq_addr       : std_logic_vector(BUS_ADDR_WIDTH-1 downto 0);
  signal Join_ss_inst_ss_net_profit_bus_rreq_len        : std_logic_vector(BUS_LEN_WIDTH-1 downto 0);
  signal Join_ss_inst_ss_net_profit_bus_rdat_valid      : std_logic;
  signal Join_ss_inst_ss_net_profit_bus_rdat_ready      : std_logic;
  signal Join_ss_inst_ss_net_profit_bus_rdat_data       : std_logic_vector(BUS_DATA_WIDTH-1 downto 0);
  signal Join_ss_inst_ss_net_profit_bus_rdat_last       : std_logic;

  signal Join_ss_inst_ss_net_profit_cmd_valid           : std_logic;
  signal Join_ss_inst_ss_net_profit_cmd_ready           : std_logic;
  signal Join_ss_inst_ss_net_profit_cmd_firstIdx        : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal Join_ss_inst_ss_net_profit_cmd_lastIdx         : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal Join_ss_inst_ss_net_profit_cmd_ctrl            : std_logic_vector(BUS_ADDR_WIDTH-1 downto 0);
  signal Join_ss_inst_ss_net_profit_cmd_tag             : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal Join_ss_inst_ss_net_profit_unl_valid           : std_logic;
  signal Join_ss_inst_ss_net_profit_unl_ready           : std_logic;
  signal Join_ss_inst_ss_net_profit_unl_tag             : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal RDAW64DW512LW8BS1BM16_inst_mst_rreq_valid      : std_logic;
  signal RDAW64DW512LW8BS1BM16_inst_mst_rreq_ready      : std_logic;
  signal RDAW64DW512LW8BS1BM16_inst_mst_rreq_addr       : std_logic_vector(BUS_ADDR_WIDTH-1 downto 0);
  signal RDAW64DW512LW8BS1BM16_inst_mst_rreq_len        : std_logic_vector(BUS_LEN_WIDTH-1 downto 0);
  signal RDAW64DW512LW8BS1BM16_inst_mst_rdat_valid      : std_logic;
  signal RDAW64DW512LW8BS1BM16_inst_mst_rdat_ready      : std_logic;
  signal RDAW64DW512LW8BS1BM16_inst_mst_rdat_data       : std_logic_vector(BUS_DATA_WIDTH-1 downto 0);
  signal RDAW64DW512LW8BS1BM16_inst_mst_rdat_last       : std_logic;

  signal RDAW64DW512LW8BS1BM16_inst_bsv_rreq_valid : std_logic_vector(6 downto 0);
  signal RDAW64DW512LW8BS1BM16_inst_bsv_rreq_ready : std_logic_vector(6 downto 0);
  signal RDAW64DW512LW8BS1BM16_inst_bsv_rreq_addr  : std_logic_vector(7*BUS_ADDR_WIDTH-1 downto 0);
  signal RDAW64DW512LW8BS1BM16_inst_bsv_rreq_len   : std_logic_vector(7*BUS_LEN_WIDTH-1 downto 0);
  signal RDAW64DW512LW8BS1BM16_inst_bsv_rdat_valid : std_logic_vector(6 downto 0);
  signal RDAW64DW512LW8BS1BM16_inst_bsv_rdat_ready : std_logic_vector(6 downto 0);
  signal RDAW64DW512LW8BS1BM16_inst_bsv_rdat_data  : std_logic_vector(7*BUS_DATA_WIDTH-1 downto 0);
  signal RDAW64DW512LW8BS1BM16_inst_bsv_rdat_last  : std_logic_vector(6 downto 0);

begin
  Join_Nucleus_inst : Join_Nucleus
    generic map (
      INDEX_WIDTH                    => INDEX_WIDTH,
      TAG_WIDTH                      => TAG_WIDTH,
      SS_SOLD_DATE_SK_BUS_ADDR_WIDTH => BUS_ADDR_WIDTH,
      SS_CDEMO_SK_BUS_ADDR_WIDTH     => BUS_ADDR_WIDTH,
      SS_ADDR_SK_BUS_ADDR_WIDTH      => BUS_ADDR_WIDTH,
      SS_STORE_SK_BUS_ADDR_WIDTH     => BUS_ADDR_WIDTH,
      SS_QUANTITY_BUS_ADDR_WIDTH     => BUS_ADDR_WIDTH,
      SS_SALES_PRICE_BUS_ADDR_WIDTH  => BUS_ADDR_WIDTH,
      SS_NET_PROFIT_BUS_ADDR_WIDTH   => BUS_ADDR_WIDTH
    )
    port map (
      kcd_clk                      => kcd_clk,
      kcd_reset                    => kcd_reset,
      mmio_awvalid                 => Join_Nucleus_inst_mmio_awvalid,
      mmio_awready                 => Join_Nucleus_inst_mmio_awready,
      mmio_awaddr                  => Join_Nucleus_inst_mmio_awaddr,
      mmio_wvalid                  => Join_Nucleus_inst_mmio_wvalid,
      mmio_wready                  => Join_Nucleus_inst_mmio_wready,
      mmio_wdata                   => Join_Nucleus_inst_mmio_wdata,
      mmio_wstrb                   => Join_Nucleus_inst_mmio_wstrb,
      mmio_bvalid                  => Join_Nucleus_inst_mmio_bvalid,
      mmio_bready                  => Join_Nucleus_inst_mmio_bready,
      mmio_bresp                   => Join_Nucleus_inst_mmio_bresp,
      mmio_arvalid                 => Join_Nucleus_inst_mmio_arvalid,
      mmio_arready                 => Join_Nucleus_inst_mmio_arready,
      mmio_araddr                  => Join_Nucleus_inst_mmio_araddr,
      mmio_rvalid                  => Join_Nucleus_inst_mmio_rvalid,
      mmio_rready                  => Join_Nucleus_inst_mmio_rready,
      mmio_rdata                   => Join_Nucleus_inst_mmio_rdata,
      mmio_rresp                   => Join_Nucleus_inst_mmio_rresp,
      ss_sold_date_sk_valid        => Join_Nucleus_inst_ss_sold_date_sk_valid,
      ss_sold_date_sk_ready        => Join_Nucleus_inst_ss_sold_date_sk_ready,
      ss_sold_date_sk_dvalid       => Join_Nucleus_inst_ss_sold_date_sk_dvalid,
      ss_sold_date_sk_last         => Join_Nucleus_inst_ss_sold_date_sk_last,
      ss_sold_date_sk              => Join_Nucleus_inst_ss_sold_date_sk,
      ss_cdemo_sk_valid            => Join_Nucleus_inst_ss_cdemo_sk_valid,
      ss_cdemo_sk_ready            => Join_Nucleus_inst_ss_cdemo_sk_ready,
      ss_cdemo_sk_dvalid           => Join_Nucleus_inst_ss_cdemo_sk_dvalid,
      ss_cdemo_sk_last             => Join_Nucleus_inst_ss_cdemo_sk_last,
      ss_cdemo_sk                  => Join_Nucleus_inst_ss_cdemo_sk,
      ss_addr_sk_valid             => Join_Nucleus_inst_ss_addr_sk_valid,
      ss_addr_sk_ready             => Join_Nucleus_inst_ss_addr_sk_ready,
      ss_addr_sk_dvalid            => Join_Nucleus_inst_ss_addr_sk_dvalid,
      ss_addr_sk_last              => Join_Nucleus_inst_ss_addr_sk_last,
      ss_addr_sk                   => Join_Nucleus_inst_ss_addr_sk,
      ss_store_sk_valid            => Join_Nucleus_inst_ss_store_sk_valid,
      ss_store_sk_ready            => Join_Nucleus_inst_ss_store_sk_ready,
      ss_store_sk_dvalid           => Join_Nucleus_inst_ss_store_sk_dvalid,
      ss_store_sk_last             => Join_Nucleus_inst_ss_store_sk_last,
      ss_store_sk                  => Join_Nucleus_inst_ss_store_sk,
      ss_quantity_valid            => Join_Nucleus_inst_ss_quantity_valid,
      ss_quantity_ready            => Join_Nucleus_inst_ss_quantity_ready,
      ss_quantity_dvalid           => Join_Nucleus_inst_ss_quantity_dvalid,
      ss_quantity_last             => Join_Nucleus_inst_ss_quantity_last,
      ss_quantity                  => Join_Nucleus_inst_ss_quantity,
      ss_sales_price_valid         => Join_Nucleus_inst_ss_sales_price_valid,
      ss_sales_price_ready         => Join_Nucleus_inst_ss_sales_price_ready,
      ss_sales_price_dvalid        => Join_Nucleus_inst_ss_sales_price_dvalid,
      ss_sales_price_last          => Join_Nucleus_inst_ss_sales_price_last,
      ss_sales_price               => Join_Nucleus_inst_ss_sales_price,
      ss_net_profit_valid          => Join_Nucleus_inst_ss_net_profit_valid,
      ss_net_profit_ready          => Join_Nucleus_inst_ss_net_profit_ready,
      ss_net_profit_dvalid         => Join_Nucleus_inst_ss_net_profit_dvalid,
      ss_net_profit_last           => Join_Nucleus_inst_ss_net_profit_last,
      ss_net_profit                => Join_Nucleus_inst_ss_net_profit,
      ss_sold_date_sk_unl_valid    => Join_Nucleus_inst_ss_sold_date_sk_unl_valid,
      ss_sold_date_sk_unl_ready    => Join_Nucleus_inst_ss_sold_date_sk_unl_ready,
      ss_sold_date_sk_unl_tag      => Join_Nucleus_inst_ss_sold_date_sk_unl_tag,
      ss_cdemo_sk_unl_valid        => Join_Nucleus_inst_ss_cdemo_sk_unl_valid,
      ss_cdemo_sk_unl_ready        => Join_Nucleus_inst_ss_cdemo_sk_unl_ready,
      ss_cdemo_sk_unl_tag          => Join_Nucleus_inst_ss_cdemo_sk_unl_tag,
      ss_addr_sk_unl_valid         => Join_Nucleus_inst_ss_addr_sk_unl_valid,
      ss_addr_sk_unl_ready         => Join_Nucleus_inst_ss_addr_sk_unl_ready,
      ss_addr_sk_unl_tag           => Join_Nucleus_inst_ss_addr_sk_unl_tag,
      ss_store_sk_unl_valid        => Join_Nucleus_inst_ss_store_sk_unl_valid,
      ss_store_sk_unl_ready        => Join_Nucleus_inst_ss_store_sk_unl_ready,
      ss_store_sk_unl_tag          => Join_Nucleus_inst_ss_store_sk_unl_tag,
      ss_quantity_unl_valid        => Join_Nucleus_inst_ss_quantity_unl_valid,
      ss_quantity_unl_ready        => Join_Nucleus_inst_ss_quantity_unl_ready,
      ss_quantity_unl_tag          => Join_Nucleus_inst_ss_quantity_unl_tag,
      ss_sales_price_unl_valid     => Join_Nucleus_inst_ss_sales_price_unl_valid,
      ss_sales_price_unl_ready     => Join_Nucleus_inst_ss_sales_price_unl_ready,
      ss_sales_price_unl_tag       => Join_Nucleus_inst_ss_sales_price_unl_tag,
      ss_net_profit_unl_valid      => Join_Nucleus_inst_ss_net_profit_unl_valid,
      ss_net_profit_unl_ready      => Join_Nucleus_inst_ss_net_profit_unl_ready,
      ss_net_profit_unl_tag        => Join_Nucleus_inst_ss_net_profit_unl_tag,
      ss_sold_date_sk_cmd_valid    => Join_Nucleus_inst_ss_sold_date_sk_cmd_valid,
      ss_sold_date_sk_cmd_ready    => Join_Nucleus_inst_ss_sold_date_sk_cmd_ready,
      ss_sold_date_sk_cmd_firstIdx => Join_Nucleus_inst_ss_sold_date_sk_cmd_firstIdx,
      ss_sold_date_sk_cmd_lastIdx  => Join_Nucleus_inst_ss_sold_date_sk_cmd_lastIdx,
      ss_sold_date_sk_cmd_ctrl     => Join_Nucleus_inst_ss_sold_date_sk_cmd_ctrl,
      ss_sold_date_sk_cmd_tag      => Join_Nucleus_inst_ss_sold_date_sk_cmd_tag,
      ss_cdemo_sk_cmd_valid        => Join_Nucleus_inst_ss_cdemo_sk_cmd_valid,
      ss_cdemo_sk_cmd_ready        => Join_Nucleus_inst_ss_cdemo_sk_cmd_ready,
      ss_cdemo_sk_cmd_firstIdx     => Join_Nucleus_inst_ss_cdemo_sk_cmd_firstIdx,
      ss_cdemo_sk_cmd_lastIdx      => Join_Nucleus_inst_ss_cdemo_sk_cmd_lastIdx,
      ss_cdemo_sk_cmd_ctrl         => Join_Nucleus_inst_ss_cdemo_sk_cmd_ctrl,
      ss_cdemo_sk_cmd_tag          => Join_Nucleus_inst_ss_cdemo_sk_cmd_tag,
      ss_addr_sk_cmd_valid         => Join_Nucleus_inst_ss_addr_sk_cmd_valid,
      ss_addr_sk_cmd_ready         => Join_Nucleus_inst_ss_addr_sk_cmd_ready,
      ss_addr_sk_cmd_firstIdx      => Join_Nucleus_inst_ss_addr_sk_cmd_firstIdx,
      ss_addr_sk_cmd_lastIdx       => Join_Nucleus_inst_ss_addr_sk_cmd_lastIdx,
      ss_addr_sk_cmd_ctrl          => Join_Nucleus_inst_ss_addr_sk_cmd_ctrl,
      ss_addr_sk_cmd_tag           => Join_Nucleus_inst_ss_addr_sk_cmd_tag,
      ss_store_sk_cmd_valid        => Join_Nucleus_inst_ss_store_sk_cmd_valid,
      ss_store_sk_cmd_ready        => Join_Nucleus_inst_ss_store_sk_cmd_ready,
      ss_store_sk_cmd_firstIdx     => Join_Nucleus_inst_ss_store_sk_cmd_firstIdx,
      ss_store_sk_cmd_lastIdx      => Join_Nucleus_inst_ss_store_sk_cmd_lastIdx,
      ss_store_sk_cmd_ctrl         => Join_Nucleus_inst_ss_store_sk_cmd_ctrl,
      ss_store_sk_cmd_tag          => Join_Nucleus_inst_ss_store_sk_cmd_tag,
      ss_quantity_cmd_valid        => Join_Nucleus_inst_ss_quantity_cmd_valid,
      ss_quantity_cmd_ready        => Join_Nucleus_inst_ss_quantity_cmd_ready,
      ss_quantity_cmd_firstIdx     => Join_Nucleus_inst_ss_quantity_cmd_firstIdx,
      ss_quantity_cmd_lastIdx      => Join_Nucleus_inst_ss_quantity_cmd_lastIdx,
      ss_quantity_cmd_ctrl         => Join_Nucleus_inst_ss_quantity_cmd_ctrl,
      ss_quantity_cmd_tag          => Join_Nucleus_inst_ss_quantity_cmd_tag,
      ss_sales_price_cmd_valid     => Join_Nucleus_inst_ss_sales_price_cmd_valid,
      ss_sales_price_cmd_ready     => Join_Nucleus_inst_ss_sales_price_cmd_ready,
      ss_sales_price_cmd_firstIdx  => Join_Nucleus_inst_ss_sales_price_cmd_firstIdx,
      ss_sales_price_cmd_lastIdx   => Join_Nucleus_inst_ss_sales_price_cmd_lastIdx,
      ss_sales_price_cmd_ctrl      => Join_Nucleus_inst_ss_sales_price_cmd_ctrl,
      ss_sales_price_cmd_tag       => Join_Nucleus_inst_ss_sales_price_cmd_tag,
      ss_net_profit_cmd_valid      => Join_Nucleus_inst_ss_net_profit_cmd_valid,
      ss_net_profit_cmd_ready      => Join_Nucleus_inst_ss_net_profit_cmd_ready,
      ss_net_profit_cmd_firstIdx   => Join_Nucleus_inst_ss_net_profit_cmd_firstIdx,
      ss_net_profit_cmd_lastIdx    => Join_Nucleus_inst_ss_net_profit_cmd_lastIdx,
      ss_net_profit_cmd_ctrl       => Join_Nucleus_inst_ss_net_profit_cmd_ctrl,
      ss_net_profit_cmd_tag        => Join_Nucleus_inst_ss_net_profit_cmd_tag
    );

  Join_ss_inst : Join_ss
    generic map (
      INDEX_WIDTH                        => INDEX_WIDTH,
      TAG_WIDTH                          => TAG_WIDTH,
      SS_SOLD_DATE_SK_BUS_ADDR_WIDTH     => BUS_ADDR_WIDTH,
      SS_SOLD_DATE_SK_BUS_DATA_WIDTH     => BUS_DATA_WIDTH,
      SS_SOLD_DATE_SK_BUS_LEN_WIDTH      => BUS_LEN_WIDTH,
      SS_SOLD_DATE_SK_BUS_BURST_STEP_LEN => BUS_BURST_STEP_LEN,
      SS_SOLD_DATE_SK_BUS_BURST_MAX_LEN  => BUS_BURST_MAX_LEN,
      SS_CDEMO_SK_BUS_ADDR_WIDTH         => BUS_ADDR_WIDTH,
      SS_CDEMO_SK_BUS_DATA_WIDTH         => BUS_DATA_WIDTH,
      SS_CDEMO_SK_BUS_LEN_WIDTH          => BUS_LEN_WIDTH,
      SS_CDEMO_SK_BUS_BURST_STEP_LEN     => BUS_BURST_STEP_LEN,
      SS_CDEMO_SK_BUS_BURST_MAX_LEN      => BUS_BURST_MAX_LEN,
      SS_ADDR_SK_BUS_ADDR_WIDTH          => BUS_ADDR_WIDTH,
      SS_ADDR_SK_BUS_DATA_WIDTH          => BUS_DATA_WIDTH,
      SS_ADDR_SK_BUS_LEN_WIDTH           => BUS_LEN_WIDTH,
      SS_ADDR_SK_BUS_BURST_STEP_LEN      => BUS_BURST_STEP_LEN,
      SS_ADDR_SK_BUS_BURST_MAX_LEN       => BUS_BURST_MAX_LEN,
      SS_STORE_SK_BUS_ADDR_WIDTH         => BUS_ADDR_WIDTH,
      SS_STORE_SK_BUS_DATA_WIDTH         => BUS_DATA_WIDTH,
      SS_STORE_SK_BUS_LEN_WIDTH          => BUS_LEN_WIDTH,
      SS_STORE_SK_BUS_BURST_STEP_LEN     => BUS_BURST_STEP_LEN,
      SS_STORE_SK_BUS_BURST_MAX_LEN      => BUS_BURST_MAX_LEN,
      SS_QUANTITY_BUS_ADDR_WIDTH         => BUS_ADDR_WIDTH,
      SS_QUANTITY_BUS_DATA_WIDTH         => BUS_DATA_WIDTH,
      SS_QUANTITY_BUS_LEN_WIDTH          => BUS_LEN_WIDTH,
      SS_QUANTITY_BUS_BURST_STEP_LEN     => BUS_BURST_STEP_LEN,
      SS_QUANTITY_BUS_BURST_MAX_LEN      => BUS_BURST_MAX_LEN,
      SS_SALES_PRICE_BUS_ADDR_WIDTH      => BUS_ADDR_WIDTH,
      SS_SALES_PRICE_BUS_DATA_WIDTH      => BUS_DATA_WIDTH,
      SS_SALES_PRICE_BUS_LEN_WIDTH       => BUS_LEN_WIDTH,
      SS_SALES_PRICE_BUS_BURST_STEP_LEN  => BUS_BURST_STEP_LEN,
      SS_SALES_PRICE_BUS_BURST_MAX_LEN   => BUS_BURST_MAX_LEN,
      SS_NET_PROFIT_BUS_ADDR_WIDTH       => BUS_ADDR_WIDTH,
      SS_NET_PROFIT_BUS_DATA_WIDTH       => BUS_DATA_WIDTH,
      SS_NET_PROFIT_BUS_LEN_WIDTH        => BUS_LEN_WIDTH,
      SS_NET_PROFIT_BUS_BURST_STEP_LEN   => BUS_BURST_STEP_LEN,
      SS_NET_PROFIT_BUS_BURST_MAX_LEN    => BUS_BURST_MAX_LEN
    )
    port map (
      bcd_clk                        => bcd_clk,
      bcd_reset                      => bcd_reset,
      kcd_clk                        => kcd_clk,
      kcd_reset                      => kcd_reset,
      ss_sold_date_sk_valid          => Join_ss_inst_ss_sold_date_sk_valid,
      ss_sold_date_sk_ready          => Join_ss_inst_ss_sold_date_sk_ready,
      ss_sold_date_sk_dvalid         => Join_ss_inst_ss_sold_date_sk_dvalid,
      ss_sold_date_sk_last           => Join_ss_inst_ss_sold_date_sk_last,
      ss_sold_date_sk                => Join_ss_inst_ss_sold_date_sk,
      ss_sold_date_sk_bus_rreq_valid => Join_ss_inst_ss_sold_date_sk_bus_rreq_valid,
      ss_sold_date_sk_bus_rreq_ready => Join_ss_inst_ss_sold_date_sk_bus_rreq_ready,
      ss_sold_date_sk_bus_rreq_addr  => Join_ss_inst_ss_sold_date_sk_bus_rreq_addr,
      ss_sold_date_sk_bus_rreq_len   => Join_ss_inst_ss_sold_date_sk_bus_rreq_len,
      ss_sold_date_sk_bus_rdat_valid => Join_ss_inst_ss_sold_date_sk_bus_rdat_valid,
      ss_sold_date_sk_bus_rdat_ready => Join_ss_inst_ss_sold_date_sk_bus_rdat_ready,
      ss_sold_date_sk_bus_rdat_data  => Join_ss_inst_ss_sold_date_sk_bus_rdat_data,
      ss_sold_date_sk_bus_rdat_last  => Join_ss_inst_ss_sold_date_sk_bus_rdat_last,
      ss_sold_date_sk_cmd_valid      => Join_ss_inst_ss_sold_date_sk_cmd_valid,
      ss_sold_date_sk_cmd_ready      => Join_ss_inst_ss_sold_date_sk_cmd_ready,
      ss_sold_date_sk_cmd_firstIdx   => Join_ss_inst_ss_sold_date_sk_cmd_firstIdx,
      ss_sold_date_sk_cmd_lastIdx    => Join_ss_inst_ss_sold_date_sk_cmd_lastIdx,
      ss_sold_date_sk_cmd_ctrl       => Join_ss_inst_ss_sold_date_sk_cmd_ctrl,
      ss_sold_date_sk_cmd_tag        => Join_ss_inst_ss_sold_date_sk_cmd_tag,
      ss_sold_date_sk_unl_valid      => Join_ss_inst_ss_sold_date_sk_unl_valid,
      ss_sold_date_sk_unl_ready      => Join_ss_inst_ss_sold_date_sk_unl_ready,
      ss_sold_date_sk_unl_tag        => Join_ss_inst_ss_sold_date_sk_unl_tag,
      ss_cdemo_sk_valid              => Join_ss_inst_ss_cdemo_sk_valid,
      ss_cdemo_sk_ready              => Join_ss_inst_ss_cdemo_sk_ready,
      ss_cdemo_sk_dvalid             => Join_ss_inst_ss_cdemo_sk_dvalid,
      ss_cdemo_sk_last               => Join_ss_inst_ss_cdemo_sk_last,
      ss_cdemo_sk                    => Join_ss_inst_ss_cdemo_sk,
      ss_cdemo_sk_bus_rreq_valid     => Join_ss_inst_ss_cdemo_sk_bus_rreq_valid,
      ss_cdemo_sk_bus_rreq_ready     => Join_ss_inst_ss_cdemo_sk_bus_rreq_ready,
      ss_cdemo_sk_bus_rreq_addr      => Join_ss_inst_ss_cdemo_sk_bus_rreq_addr,
      ss_cdemo_sk_bus_rreq_len       => Join_ss_inst_ss_cdemo_sk_bus_rreq_len,
      ss_cdemo_sk_bus_rdat_valid     => Join_ss_inst_ss_cdemo_sk_bus_rdat_valid,
      ss_cdemo_sk_bus_rdat_ready     => Join_ss_inst_ss_cdemo_sk_bus_rdat_ready,
      ss_cdemo_sk_bus_rdat_data      => Join_ss_inst_ss_cdemo_sk_bus_rdat_data,
      ss_cdemo_sk_bus_rdat_last      => Join_ss_inst_ss_cdemo_sk_bus_rdat_last,
      ss_cdemo_sk_cmd_valid          => Join_ss_inst_ss_cdemo_sk_cmd_valid,
      ss_cdemo_sk_cmd_ready          => Join_ss_inst_ss_cdemo_sk_cmd_ready,
      ss_cdemo_sk_cmd_firstIdx       => Join_ss_inst_ss_cdemo_sk_cmd_firstIdx,
      ss_cdemo_sk_cmd_lastIdx        => Join_ss_inst_ss_cdemo_sk_cmd_lastIdx,
      ss_cdemo_sk_cmd_ctrl           => Join_ss_inst_ss_cdemo_sk_cmd_ctrl,
      ss_cdemo_sk_cmd_tag            => Join_ss_inst_ss_cdemo_sk_cmd_tag,
      ss_cdemo_sk_unl_valid          => Join_ss_inst_ss_cdemo_sk_unl_valid,
      ss_cdemo_sk_unl_ready          => Join_ss_inst_ss_cdemo_sk_unl_ready,
      ss_cdemo_sk_unl_tag            => Join_ss_inst_ss_cdemo_sk_unl_tag,
      ss_addr_sk_valid               => Join_ss_inst_ss_addr_sk_valid,
      ss_addr_sk_ready               => Join_ss_inst_ss_addr_sk_ready,
      ss_addr_sk_dvalid              => Join_ss_inst_ss_addr_sk_dvalid,
      ss_addr_sk_last                => Join_ss_inst_ss_addr_sk_last,
      ss_addr_sk                     => Join_ss_inst_ss_addr_sk,
      ss_addr_sk_bus_rreq_valid      => Join_ss_inst_ss_addr_sk_bus_rreq_valid,
      ss_addr_sk_bus_rreq_ready      => Join_ss_inst_ss_addr_sk_bus_rreq_ready,
      ss_addr_sk_bus_rreq_addr       => Join_ss_inst_ss_addr_sk_bus_rreq_addr,
      ss_addr_sk_bus_rreq_len        => Join_ss_inst_ss_addr_sk_bus_rreq_len,
      ss_addr_sk_bus_rdat_valid      => Join_ss_inst_ss_addr_sk_bus_rdat_valid,
      ss_addr_sk_bus_rdat_ready      => Join_ss_inst_ss_addr_sk_bus_rdat_ready,
      ss_addr_sk_bus_rdat_data       => Join_ss_inst_ss_addr_sk_bus_rdat_data,
      ss_addr_sk_bus_rdat_last       => Join_ss_inst_ss_addr_sk_bus_rdat_last,
      ss_addr_sk_cmd_valid           => Join_ss_inst_ss_addr_sk_cmd_valid,
      ss_addr_sk_cmd_ready           => Join_ss_inst_ss_addr_sk_cmd_ready,
      ss_addr_sk_cmd_firstIdx        => Join_ss_inst_ss_addr_sk_cmd_firstIdx,
      ss_addr_sk_cmd_lastIdx         => Join_ss_inst_ss_addr_sk_cmd_lastIdx,
      ss_addr_sk_cmd_ctrl            => Join_ss_inst_ss_addr_sk_cmd_ctrl,
      ss_addr_sk_cmd_tag             => Join_ss_inst_ss_addr_sk_cmd_tag,
      ss_addr_sk_unl_valid           => Join_ss_inst_ss_addr_sk_unl_valid,
      ss_addr_sk_unl_ready           => Join_ss_inst_ss_addr_sk_unl_ready,
      ss_addr_sk_unl_tag             => Join_ss_inst_ss_addr_sk_unl_tag,
      ss_store_sk_valid              => Join_ss_inst_ss_store_sk_valid,
      ss_store_sk_ready              => Join_ss_inst_ss_store_sk_ready,
      ss_store_sk_dvalid             => Join_ss_inst_ss_store_sk_dvalid,
      ss_store_sk_last               => Join_ss_inst_ss_store_sk_last,
      ss_store_sk                    => Join_ss_inst_ss_store_sk,
      ss_store_sk_bus_rreq_valid     => Join_ss_inst_ss_store_sk_bus_rreq_valid,
      ss_store_sk_bus_rreq_ready     => Join_ss_inst_ss_store_sk_bus_rreq_ready,
      ss_store_sk_bus_rreq_addr      => Join_ss_inst_ss_store_sk_bus_rreq_addr,
      ss_store_sk_bus_rreq_len       => Join_ss_inst_ss_store_sk_bus_rreq_len,
      ss_store_sk_bus_rdat_valid     => Join_ss_inst_ss_store_sk_bus_rdat_valid,
      ss_store_sk_bus_rdat_ready     => Join_ss_inst_ss_store_sk_bus_rdat_ready,
      ss_store_sk_bus_rdat_data      => Join_ss_inst_ss_store_sk_bus_rdat_data,
      ss_store_sk_bus_rdat_last      => Join_ss_inst_ss_store_sk_bus_rdat_last,
      ss_store_sk_cmd_valid          => Join_ss_inst_ss_store_sk_cmd_valid,
      ss_store_sk_cmd_ready          => Join_ss_inst_ss_store_sk_cmd_ready,
      ss_store_sk_cmd_firstIdx       => Join_ss_inst_ss_store_sk_cmd_firstIdx,
      ss_store_sk_cmd_lastIdx        => Join_ss_inst_ss_store_sk_cmd_lastIdx,
      ss_store_sk_cmd_ctrl           => Join_ss_inst_ss_store_sk_cmd_ctrl,
      ss_store_sk_cmd_tag            => Join_ss_inst_ss_store_sk_cmd_tag,
      ss_store_sk_unl_valid          => Join_ss_inst_ss_store_sk_unl_valid,
      ss_store_sk_unl_ready          => Join_ss_inst_ss_store_sk_unl_ready,
      ss_store_sk_unl_tag            => Join_ss_inst_ss_store_sk_unl_tag,
      ss_quantity_valid              => Join_ss_inst_ss_quantity_valid,
      ss_quantity_ready              => Join_ss_inst_ss_quantity_ready,
      ss_quantity_dvalid             => Join_ss_inst_ss_quantity_dvalid,
      ss_quantity_last               => Join_ss_inst_ss_quantity_last,
      ss_quantity                    => Join_ss_inst_ss_quantity,
      ss_quantity_bus_rreq_valid     => Join_ss_inst_ss_quantity_bus_rreq_valid,
      ss_quantity_bus_rreq_ready     => Join_ss_inst_ss_quantity_bus_rreq_ready,
      ss_quantity_bus_rreq_addr      => Join_ss_inst_ss_quantity_bus_rreq_addr,
      ss_quantity_bus_rreq_len       => Join_ss_inst_ss_quantity_bus_rreq_len,
      ss_quantity_bus_rdat_valid     => Join_ss_inst_ss_quantity_bus_rdat_valid,
      ss_quantity_bus_rdat_ready     => Join_ss_inst_ss_quantity_bus_rdat_ready,
      ss_quantity_bus_rdat_data      => Join_ss_inst_ss_quantity_bus_rdat_data,
      ss_quantity_bus_rdat_last      => Join_ss_inst_ss_quantity_bus_rdat_last,
      ss_quantity_cmd_valid          => Join_ss_inst_ss_quantity_cmd_valid,
      ss_quantity_cmd_ready          => Join_ss_inst_ss_quantity_cmd_ready,
      ss_quantity_cmd_firstIdx       => Join_ss_inst_ss_quantity_cmd_firstIdx,
      ss_quantity_cmd_lastIdx        => Join_ss_inst_ss_quantity_cmd_lastIdx,
      ss_quantity_cmd_ctrl           => Join_ss_inst_ss_quantity_cmd_ctrl,
      ss_quantity_cmd_tag            => Join_ss_inst_ss_quantity_cmd_tag,
      ss_quantity_unl_valid          => Join_ss_inst_ss_quantity_unl_valid,
      ss_quantity_unl_ready          => Join_ss_inst_ss_quantity_unl_ready,
      ss_quantity_unl_tag            => Join_ss_inst_ss_quantity_unl_tag,
      ss_sales_price_valid           => Join_ss_inst_ss_sales_price_valid,
      ss_sales_price_ready           => Join_ss_inst_ss_sales_price_ready,
      ss_sales_price_dvalid          => Join_ss_inst_ss_sales_price_dvalid,
      ss_sales_price_last            => Join_ss_inst_ss_sales_price_last,
      ss_sales_price                 => Join_ss_inst_ss_sales_price,
      ss_sales_price_bus_rreq_valid  => Join_ss_inst_ss_sales_price_bus_rreq_valid,
      ss_sales_price_bus_rreq_ready  => Join_ss_inst_ss_sales_price_bus_rreq_ready,
      ss_sales_price_bus_rreq_addr   => Join_ss_inst_ss_sales_price_bus_rreq_addr,
      ss_sales_price_bus_rreq_len    => Join_ss_inst_ss_sales_price_bus_rreq_len,
      ss_sales_price_bus_rdat_valid  => Join_ss_inst_ss_sales_price_bus_rdat_valid,
      ss_sales_price_bus_rdat_ready  => Join_ss_inst_ss_sales_price_bus_rdat_ready,
      ss_sales_price_bus_rdat_data   => Join_ss_inst_ss_sales_price_bus_rdat_data,
      ss_sales_price_bus_rdat_last   => Join_ss_inst_ss_sales_price_bus_rdat_last,
      ss_sales_price_cmd_valid       => Join_ss_inst_ss_sales_price_cmd_valid,
      ss_sales_price_cmd_ready       => Join_ss_inst_ss_sales_price_cmd_ready,
      ss_sales_price_cmd_firstIdx    => Join_ss_inst_ss_sales_price_cmd_firstIdx,
      ss_sales_price_cmd_lastIdx     => Join_ss_inst_ss_sales_price_cmd_lastIdx,
      ss_sales_price_cmd_ctrl        => Join_ss_inst_ss_sales_price_cmd_ctrl,
      ss_sales_price_cmd_tag         => Join_ss_inst_ss_sales_price_cmd_tag,
      ss_sales_price_unl_valid       => Join_ss_inst_ss_sales_price_unl_valid,
      ss_sales_price_unl_ready       => Join_ss_inst_ss_sales_price_unl_ready,
      ss_sales_price_unl_tag         => Join_ss_inst_ss_sales_price_unl_tag,
      ss_net_profit_valid            => Join_ss_inst_ss_net_profit_valid,
      ss_net_profit_ready            => Join_ss_inst_ss_net_profit_ready,
      ss_net_profit_dvalid           => Join_ss_inst_ss_net_profit_dvalid,
      ss_net_profit_last             => Join_ss_inst_ss_net_profit_last,
      ss_net_profit                  => Join_ss_inst_ss_net_profit,
      ss_net_profit_bus_rreq_valid   => Join_ss_inst_ss_net_profit_bus_rreq_valid,
      ss_net_profit_bus_rreq_ready   => Join_ss_inst_ss_net_profit_bus_rreq_ready,
      ss_net_profit_bus_rreq_addr    => Join_ss_inst_ss_net_profit_bus_rreq_addr,
      ss_net_profit_bus_rreq_len     => Join_ss_inst_ss_net_profit_bus_rreq_len,
      ss_net_profit_bus_rdat_valid   => Join_ss_inst_ss_net_profit_bus_rdat_valid,
      ss_net_profit_bus_rdat_ready   => Join_ss_inst_ss_net_profit_bus_rdat_ready,
      ss_net_profit_bus_rdat_data    => Join_ss_inst_ss_net_profit_bus_rdat_data,
      ss_net_profit_bus_rdat_last    => Join_ss_inst_ss_net_profit_bus_rdat_last,
      ss_net_profit_cmd_valid        => Join_ss_inst_ss_net_profit_cmd_valid,
      ss_net_profit_cmd_ready        => Join_ss_inst_ss_net_profit_cmd_ready,
      ss_net_profit_cmd_firstIdx     => Join_ss_inst_ss_net_profit_cmd_firstIdx,
      ss_net_profit_cmd_lastIdx      => Join_ss_inst_ss_net_profit_cmd_lastIdx,
      ss_net_profit_cmd_ctrl         => Join_ss_inst_ss_net_profit_cmd_ctrl,
      ss_net_profit_cmd_tag          => Join_ss_inst_ss_net_profit_cmd_tag,
      ss_net_profit_unl_valid        => Join_ss_inst_ss_net_profit_unl_valid,
      ss_net_profit_unl_ready        => Join_ss_inst_ss_net_profit_unl_ready,
      ss_net_profit_unl_tag          => Join_ss_inst_ss_net_profit_unl_tag
    );

  RDAW64DW512LW8BS1BM16_inst : BusReadArbiterVec
    generic map (
      BUS_ADDR_WIDTH  => BUS_ADDR_WIDTH,
      BUS_DATA_WIDTH  => BUS_DATA_WIDTH,
      BUS_LEN_WIDTH   => BUS_LEN_WIDTH,
      NUM_SLAVE_PORTS => 7,
      ARB_METHOD      => "RR-STICKY",
      MAX_OUTSTANDING => 4,
      RAM_CONFIG      => "",
      SLV_REQ_SLICES  => true,
      MST_REQ_SLICE   => true,
      MST_DAT_SLICE   => true,
      SLV_DAT_SLICES  => true
    )
    port map (
      bcd_clk        => bcd_clk,
      bcd_reset      => bcd_reset,
      mst_rreq_valid => RDAW64DW512LW8BS1BM16_inst_mst_rreq_valid,
      mst_rreq_ready => RDAW64DW512LW8BS1BM16_inst_mst_rreq_ready,
      mst_rreq_addr  => RDAW64DW512LW8BS1BM16_inst_mst_rreq_addr,
      mst_rreq_len   => RDAW64DW512LW8BS1BM16_inst_mst_rreq_len,
      mst_rdat_valid => RDAW64DW512LW8BS1BM16_inst_mst_rdat_valid,
      mst_rdat_ready => RDAW64DW512LW8BS1BM16_inst_mst_rdat_ready,
      mst_rdat_data  => RDAW64DW512LW8BS1BM16_inst_mst_rdat_data,
      mst_rdat_last  => RDAW64DW512LW8BS1BM16_inst_mst_rdat_last,
      bsv_rreq_valid => RDAW64DW512LW8BS1BM16_inst_bsv_rreq_valid,
      bsv_rreq_ready => RDAW64DW512LW8BS1BM16_inst_bsv_rreq_ready,
      bsv_rreq_len   => RDAW64DW512LW8BS1BM16_inst_bsv_rreq_len,
      bsv_rreq_addr  => RDAW64DW512LW8BS1BM16_inst_bsv_rreq_addr,
      bsv_rdat_valid => RDAW64DW512LW8BS1BM16_inst_bsv_rdat_valid,
      bsv_rdat_ready => RDAW64DW512LW8BS1BM16_inst_bsv_rdat_ready,
      bsv_rdat_last  => RDAW64DW512LW8BS1BM16_inst_bsv_rdat_last,
      bsv_rdat_data  => RDAW64DW512LW8BS1BM16_inst_bsv_rdat_data
    );

  rd_mst_rreq_valid                         <= RDAW64DW512LW8BS1BM16_inst_mst_rreq_valid;
  RDAW64DW512LW8BS1BM16_inst_mst_rreq_ready <= rd_mst_rreq_ready;
  rd_mst_rreq_addr                          <= RDAW64DW512LW8BS1BM16_inst_mst_rreq_addr;
  rd_mst_rreq_len                           <= RDAW64DW512LW8BS1BM16_inst_mst_rreq_len;
  RDAW64DW512LW8BS1BM16_inst_mst_rdat_valid <= rd_mst_rdat_valid;
  rd_mst_rdat_ready                         <= RDAW64DW512LW8BS1BM16_inst_mst_rdat_ready;
  RDAW64DW512LW8BS1BM16_inst_mst_rdat_data  <= rd_mst_rdat_data;
  RDAW64DW512LW8BS1BM16_inst_mst_rdat_last  <= rd_mst_rdat_last;

  Join_Nucleus_inst_mmio_awvalid              <= mmio_awvalid;
  mmio_awready                                <= Join_Nucleus_inst_mmio_awready;
  Join_Nucleus_inst_mmio_awaddr               <= mmio_awaddr;
  Join_Nucleus_inst_mmio_wvalid               <= mmio_wvalid;
  mmio_wready                                 <= Join_Nucleus_inst_mmio_wready;
  Join_Nucleus_inst_mmio_wdata                <= mmio_wdata;
  Join_Nucleus_inst_mmio_wstrb                <= mmio_wstrb;
  mmio_bvalid                                 <= Join_Nucleus_inst_mmio_bvalid;
  Join_Nucleus_inst_mmio_bready               <= mmio_bready;
  mmio_bresp                                  <= Join_Nucleus_inst_mmio_bresp;
  Join_Nucleus_inst_mmio_arvalid              <= mmio_arvalid;
  mmio_arready                                <= Join_Nucleus_inst_mmio_arready;
  Join_Nucleus_inst_mmio_araddr               <= mmio_araddr;
  mmio_rvalid                                 <= Join_Nucleus_inst_mmio_rvalid;
  Join_Nucleus_inst_mmio_rready               <= mmio_rready;
  mmio_rdata                                  <= Join_Nucleus_inst_mmio_rdata;
  mmio_rresp                                  <= Join_Nucleus_inst_mmio_rresp;

  Join_Nucleus_inst_ss_sold_date_sk_valid     <= Join_ss_inst_ss_sold_date_sk_valid;
  Join_ss_inst_ss_sold_date_sk_ready          <= Join_Nucleus_inst_ss_sold_date_sk_ready;
  Join_Nucleus_inst_ss_sold_date_sk_dvalid    <= Join_ss_inst_ss_sold_date_sk_dvalid;
  Join_Nucleus_inst_ss_sold_date_sk_last      <= Join_ss_inst_ss_sold_date_sk_last;
  Join_Nucleus_inst_ss_sold_date_sk           <= Join_ss_inst_ss_sold_date_sk;

  Join_Nucleus_inst_ss_cdemo_sk_valid         <= Join_ss_inst_ss_cdemo_sk_valid;
  Join_ss_inst_ss_cdemo_sk_ready              <= Join_Nucleus_inst_ss_cdemo_sk_ready;
  Join_Nucleus_inst_ss_cdemo_sk_dvalid        <= Join_ss_inst_ss_cdemo_sk_dvalid;
  Join_Nucleus_inst_ss_cdemo_sk_last          <= Join_ss_inst_ss_cdemo_sk_last;
  Join_Nucleus_inst_ss_cdemo_sk               <= Join_ss_inst_ss_cdemo_sk;

  Join_Nucleus_inst_ss_addr_sk_valid          <= Join_ss_inst_ss_addr_sk_valid;
  Join_ss_inst_ss_addr_sk_ready               <= Join_Nucleus_inst_ss_addr_sk_ready;
  Join_Nucleus_inst_ss_addr_sk_dvalid         <= Join_ss_inst_ss_addr_sk_dvalid;
  Join_Nucleus_inst_ss_addr_sk_last           <= Join_ss_inst_ss_addr_sk_last;
  Join_Nucleus_inst_ss_addr_sk                <= Join_ss_inst_ss_addr_sk;

  Join_Nucleus_inst_ss_store_sk_valid         <= Join_ss_inst_ss_store_sk_valid;
  Join_ss_inst_ss_store_sk_ready              <= Join_Nucleus_inst_ss_store_sk_ready;
  Join_Nucleus_inst_ss_store_sk_dvalid        <= Join_ss_inst_ss_store_sk_dvalid;
  Join_Nucleus_inst_ss_store_sk_last          <= Join_ss_inst_ss_store_sk_last;
  Join_Nucleus_inst_ss_store_sk               <= Join_ss_inst_ss_store_sk;

  Join_Nucleus_inst_ss_quantity_valid         <= Join_ss_inst_ss_quantity_valid;
  Join_ss_inst_ss_quantity_ready              <= Join_Nucleus_inst_ss_quantity_ready;
  Join_Nucleus_inst_ss_quantity_dvalid        <= Join_ss_inst_ss_quantity_dvalid;
  Join_Nucleus_inst_ss_quantity_last          <= Join_ss_inst_ss_quantity_last;
  Join_Nucleus_inst_ss_quantity               <= Join_ss_inst_ss_quantity;

  Join_Nucleus_inst_ss_sales_price_valid      <= Join_ss_inst_ss_sales_price_valid;
  Join_ss_inst_ss_sales_price_ready           <= Join_Nucleus_inst_ss_sales_price_ready;
  Join_Nucleus_inst_ss_sales_price_dvalid     <= Join_ss_inst_ss_sales_price_dvalid;
  Join_Nucleus_inst_ss_sales_price_last       <= Join_ss_inst_ss_sales_price_last;
  Join_Nucleus_inst_ss_sales_price            <= Join_ss_inst_ss_sales_price;

  Join_Nucleus_inst_ss_net_profit_valid       <= Join_ss_inst_ss_net_profit_valid;
  Join_ss_inst_ss_net_profit_ready            <= Join_Nucleus_inst_ss_net_profit_ready;
  Join_Nucleus_inst_ss_net_profit_dvalid      <= Join_ss_inst_ss_net_profit_dvalid;
  Join_Nucleus_inst_ss_net_profit_last        <= Join_ss_inst_ss_net_profit_last;
  Join_Nucleus_inst_ss_net_profit             <= Join_ss_inst_ss_net_profit;

  Join_Nucleus_inst_ss_sold_date_sk_unl_valid <= Join_ss_inst_ss_sold_date_sk_unl_valid;
  Join_ss_inst_ss_sold_date_sk_unl_ready      <= Join_Nucleus_inst_ss_sold_date_sk_unl_ready;
  Join_Nucleus_inst_ss_sold_date_sk_unl_tag   <= Join_ss_inst_ss_sold_date_sk_unl_tag;

  Join_Nucleus_inst_ss_cdemo_sk_unl_valid     <= Join_ss_inst_ss_cdemo_sk_unl_valid;
  Join_ss_inst_ss_cdemo_sk_unl_ready          <= Join_Nucleus_inst_ss_cdemo_sk_unl_ready;
  Join_Nucleus_inst_ss_cdemo_sk_unl_tag       <= Join_ss_inst_ss_cdemo_sk_unl_tag;

  Join_Nucleus_inst_ss_addr_sk_unl_valid      <= Join_ss_inst_ss_addr_sk_unl_valid;
  Join_ss_inst_ss_addr_sk_unl_ready           <= Join_Nucleus_inst_ss_addr_sk_unl_ready;
  Join_Nucleus_inst_ss_addr_sk_unl_tag        <= Join_ss_inst_ss_addr_sk_unl_tag;

  Join_Nucleus_inst_ss_store_sk_unl_valid     <= Join_ss_inst_ss_store_sk_unl_valid;
  Join_ss_inst_ss_store_sk_unl_ready          <= Join_Nucleus_inst_ss_store_sk_unl_ready;
  Join_Nucleus_inst_ss_store_sk_unl_tag       <= Join_ss_inst_ss_store_sk_unl_tag;

  Join_Nucleus_inst_ss_quantity_unl_valid     <= Join_ss_inst_ss_quantity_unl_valid;
  Join_ss_inst_ss_quantity_unl_ready          <= Join_Nucleus_inst_ss_quantity_unl_ready;
  Join_Nucleus_inst_ss_quantity_unl_tag       <= Join_ss_inst_ss_quantity_unl_tag;

  Join_Nucleus_inst_ss_sales_price_unl_valid  <= Join_ss_inst_ss_sales_price_unl_valid;
  Join_ss_inst_ss_sales_price_unl_ready       <= Join_Nucleus_inst_ss_sales_price_unl_ready;
  Join_Nucleus_inst_ss_sales_price_unl_tag    <= Join_ss_inst_ss_sales_price_unl_tag;

  Join_Nucleus_inst_ss_net_profit_unl_valid   <= Join_ss_inst_ss_net_profit_unl_valid;
  Join_ss_inst_ss_net_profit_unl_ready        <= Join_Nucleus_inst_ss_net_profit_unl_ready;
  Join_Nucleus_inst_ss_net_profit_unl_tag     <= Join_ss_inst_ss_net_profit_unl_tag;

  Join_ss_inst_ss_sold_date_sk_cmd_valid      <= Join_Nucleus_inst_ss_sold_date_sk_cmd_valid;
  Join_Nucleus_inst_ss_sold_date_sk_cmd_ready <= Join_ss_inst_ss_sold_date_sk_cmd_ready;
  Join_ss_inst_ss_sold_date_sk_cmd_firstIdx   <= Join_Nucleus_inst_ss_sold_date_sk_cmd_firstIdx;
  Join_ss_inst_ss_sold_date_sk_cmd_lastIdx    <= Join_Nucleus_inst_ss_sold_date_sk_cmd_lastIdx;
  Join_ss_inst_ss_sold_date_sk_cmd_ctrl       <= Join_Nucleus_inst_ss_sold_date_sk_cmd_ctrl;
  Join_ss_inst_ss_sold_date_sk_cmd_tag        <= Join_Nucleus_inst_ss_sold_date_sk_cmd_tag;

  Join_ss_inst_ss_cdemo_sk_cmd_valid          <= Join_Nucleus_inst_ss_cdemo_sk_cmd_valid;
  Join_Nucleus_inst_ss_cdemo_sk_cmd_ready     <= Join_ss_inst_ss_cdemo_sk_cmd_ready;
  Join_ss_inst_ss_cdemo_sk_cmd_firstIdx       <= Join_Nucleus_inst_ss_cdemo_sk_cmd_firstIdx;
  Join_ss_inst_ss_cdemo_sk_cmd_lastIdx        <= Join_Nucleus_inst_ss_cdemo_sk_cmd_lastIdx;
  Join_ss_inst_ss_cdemo_sk_cmd_ctrl           <= Join_Nucleus_inst_ss_cdemo_sk_cmd_ctrl;
  Join_ss_inst_ss_cdemo_sk_cmd_tag            <= Join_Nucleus_inst_ss_cdemo_sk_cmd_tag;

  Join_ss_inst_ss_addr_sk_cmd_valid           <= Join_Nucleus_inst_ss_addr_sk_cmd_valid;
  Join_Nucleus_inst_ss_addr_sk_cmd_ready      <= Join_ss_inst_ss_addr_sk_cmd_ready;
  Join_ss_inst_ss_addr_sk_cmd_firstIdx        <= Join_Nucleus_inst_ss_addr_sk_cmd_firstIdx;
  Join_ss_inst_ss_addr_sk_cmd_lastIdx         <= Join_Nucleus_inst_ss_addr_sk_cmd_lastIdx;
  Join_ss_inst_ss_addr_sk_cmd_ctrl            <= Join_Nucleus_inst_ss_addr_sk_cmd_ctrl;
  Join_ss_inst_ss_addr_sk_cmd_tag             <= Join_Nucleus_inst_ss_addr_sk_cmd_tag;

  Join_ss_inst_ss_store_sk_cmd_valid          <= Join_Nucleus_inst_ss_store_sk_cmd_valid;
  Join_Nucleus_inst_ss_store_sk_cmd_ready     <= Join_ss_inst_ss_store_sk_cmd_ready;
  Join_ss_inst_ss_store_sk_cmd_firstIdx       <= Join_Nucleus_inst_ss_store_sk_cmd_firstIdx;
  Join_ss_inst_ss_store_sk_cmd_lastIdx        <= Join_Nucleus_inst_ss_store_sk_cmd_lastIdx;
  Join_ss_inst_ss_store_sk_cmd_ctrl           <= Join_Nucleus_inst_ss_store_sk_cmd_ctrl;
  Join_ss_inst_ss_store_sk_cmd_tag            <= Join_Nucleus_inst_ss_store_sk_cmd_tag;

  Join_ss_inst_ss_quantity_cmd_valid          <= Join_Nucleus_inst_ss_quantity_cmd_valid;
  Join_Nucleus_inst_ss_quantity_cmd_ready     <= Join_ss_inst_ss_quantity_cmd_ready;
  Join_ss_inst_ss_quantity_cmd_firstIdx       <= Join_Nucleus_inst_ss_quantity_cmd_firstIdx;
  Join_ss_inst_ss_quantity_cmd_lastIdx        <= Join_Nucleus_inst_ss_quantity_cmd_lastIdx;
  Join_ss_inst_ss_quantity_cmd_ctrl           <= Join_Nucleus_inst_ss_quantity_cmd_ctrl;
  Join_ss_inst_ss_quantity_cmd_tag            <= Join_Nucleus_inst_ss_quantity_cmd_tag;

  Join_ss_inst_ss_sales_price_cmd_valid       <= Join_Nucleus_inst_ss_sales_price_cmd_valid;
  Join_Nucleus_inst_ss_sales_price_cmd_ready  <= Join_ss_inst_ss_sales_price_cmd_ready;
  Join_ss_inst_ss_sales_price_cmd_firstIdx    <= Join_Nucleus_inst_ss_sales_price_cmd_firstIdx;
  Join_ss_inst_ss_sales_price_cmd_lastIdx     <= Join_Nucleus_inst_ss_sales_price_cmd_lastIdx;
  Join_ss_inst_ss_sales_price_cmd_ctrl        <= Join_Nucleus_inst_ss_sales_price_cmd_ctrl;
  Join_ss_inst_ss_sales_price_cmd_tag         <= Join_Nucleus_inst_ss_sales_price_cmd_tag;

  Join_ss_inst_ss_net_profit_cmd_valid        <= Join_Nucleus_inst_ss_net_profit_cmd_valid;
  Join_Nucleus_inst_ss_net_profit_cmd_ready   <= Join_ss_inst_ss_net_profit_cmd_ready;
  Join_ss_inst_ss_net_profit_cmd_firstIdx     <= Join_Nucleus_inst_ss_net_profit_cmd_firstIdx;
  Join_ss_inst_ss_net_profit_cmd_lastIdx      <= Join_Nucleus_inst_ss_net_profit_cmd_lastIdx;
  Join_ss_inst_ss_net_profit_cmd_ctrl         <= Join_Nucleus_inst_ss_net_profit_cmd_ctrl;
  Join_ss_inst_ss_net_profit_cmd_tag          <= Join_Nucleus_inst_ss_net_profit_cmd_tag;

  RDAW64DW512LW8BS1BM16_inst_bsv_rreq_valid(0)                                                        <= Join_ss_inst_ss_sold_date_sk_bus_rreq_valid;
  RDAW64DW512LW8BS1BM16_inst_bsv_rreq_valid(1)                                                        <= Join_ss_inst_ss_cdemo_sk_bus_rreq_valid;
  RDAW64DW512LW8BS1BM16_inst_bsv_rreq_valid(2)                                                        <= Join_ss_inst_ss_addr_sk_bus_rreq_valid;
  RDAW64DW512LW8BS1BM16_inst_bsv_rreq_valid(3)                                                        <= Join_ss_inst_ss_store_sk_bus_rreq_valid;
  RDAW64DW512LW8BS1BM16_inst_bsv_rreq_valid(4)                                                        <= Join_ss_inst_ss_quantity_bus_rreq_valid;
  RDAW64DW512LW8BS1BM16_inst_bsv_rreq_valid(5)                                                        <= Join_ss_inst_ss_sales_price_bus_rreq_valid;
  RDAW64DW512LW8BS1BM16_inst_bsv_rreq_valid(6)                                                        <= Join_ss_inst_ss_net_profit_bus_rreq_valid;
  RDAW64DW512LW8BS1BM16_inst_bsv_rreq_len(BUS_LEN_WIDTH-1 downto 0)                                   <= Join_ss_inst_ss_sold_date_sk_bus_rreq_len;
  RDAW64DW512LW8BS1BM16_inst_bsv_rreq_len(BUS_LEN_WIDTH+BUS_LEN_WIDTH-1 downto BUS_LEN_WIDTH)         <= Join_ss_inst_ss_cdemo_sk_bus_rreq_len;
  RDAW64DW512LW8BS1BM16_inst_bsv_rreq_len(BUS_LEN_WIDTH*2+BUS_LEN_WIDTH-1 downto BUS_LEN_WIDTH*2)     <= Join_ss_inst_ss_addr_sk_bus_rreq_len;
  RDAW64DW512LW8BS1BM16_inst_bsv_rreq_len(BUS_LEN_WIDTH*3+BUS_LEN_WIDTH-1 downto BUS_LEN_WIDTH*3)     <= Join_ss_inst_ss_store_sk_bus_rreq_len;
  RDAW64DW512LW8BS1BM16_inst_bsv_rreq_len(BUS_LEN_WIDTH*4+BUS_LEN_WIDTH-1 downto BUS_LEN_WIDTH*4)     <= Join_ss_inst_ss_quantity_bus_rreq_len;
  RDAW64DW512LW8BS1BM16_inst_bsv_rreq_len(BUS_LEN_WIDTH*5+BUS_LEN_WIDTH-1 downto BUS_LEN_WIDTH*5)     <= Join_ss_inst_ss_sales_price_bus_rreq_len;
  RDAW64DW512LW8BS1BM16_inst_bsv_rreq_len(BUS_LEN_WIDTH*6+BUS_LEN_WIDTH-1 downto BUS_LEN_WIDTH*6)     <= Join_ss_inst_ss_net_profit_bus_rreq_len;
  RDAW64DW512LW8BS1BM16_inst_bsv_rreq_addr(BUS_ADDR_WIDTH-1 downto 0)                                 <= Join_ss_inst_ss_sold_date_sk_bus_rreq_addr;
  RDAW64DW512LW8BS1BM16_inst_bsv_rreq_addr(BUS_ADDR_WIDTH+BUS_ADDR_WIDTH-1 downto BUS_ADDR_WIDTH)     <= Join_ss_inst_ss_cdemo_sk_bus_rreq_addr;
  RDAW64DW512LW8BS1BM16_inst_bsv_rreq_addr(BUS_ADDR_WIDTH*2+BUS_ADDR_WIDTH-1 downto BUS_ADDR_WIDTH*2) <= Join_ss_inst_ss_addr_sk_bus_rreq_addr;
  RDAW64DW512LW8BS1BM16_inst_bsv_rreq_addr(BUS_ADDR_WIDTH*3+BUS_ADDR_WIDTH-1 downto BUS_ADDR_WIDTH*3) <= Join_ss_inst_ss_store_sk_bus_rreq_addr;
  RDAW64DW512LW8BS1BM16_inst_bsv_rreq_addr(BUS_ADDR_WIDTH*4+BUS_ADDR_WIDTH-1 downto BUS_ADDR_WIDTH*4) <= Join_ss_inst_ss_quantity_bus_rreq_addr;
  RDAW64DW512LW8BS1BM16_inst_bsv_rreq_addr(BUS_ADDR_WIDTH*5+BUS_ADDR_WIDTH-1 downto BUS_ADDR_WIDTH*5) <= Join_ss_inst_ss_sales_price_bus_rreq_addr;
  RDAW64DW512LW8BS1BM16_inst_bsv_rreq_addr(BUS_ADDR_WIDTH*6+BUS_ADDR_WIDTH-1 downto BUS_ADDR_WIDTH*6) <= Join_ss_inst_ss_net_profit_bus_rreq_addr;
  RDAW64DW512LW8BS1BM16_inst_bsv_rdat_ready(0)                                                        <= Join_ss_inst_ss_sold_date_sk_bus_rdat_ready;
  RDAW64DW512LW8BS1BM16_inst_bsv_rdat_ready(1)                                                        <= Join_ss_inst_ss_cdemo_sk_bus_rdat_ready;
  RDAW64DW512LW8BS1BM16_inst_bsv_rdat_ready(2)                                                        <= Join_ss_inst_ss_addr_sk_bus_rdat_ready;
  RDAW64DW512LW8BS1BM16_inst_bsv_rdat_ready(3)                                                        <= Join_ss_inst_ss_store_sk_bus_rdat_ready;
  RDAW64DW512LW8BS1BM16_inst_bsv_rdat_ready(4)                                                        <= Join_ss_inst_ss_quantity_bus_rdat_ready;
  RDAW64DW512LW8BS1BM16_inst_bsv_rdat_ready(5)                                                        <= Join_ss_inst_ss_sales_price_bus_rdat_ready;
  RDAW64DW512LW8BS1BM16_inst_bsv_rdat_ready(6)                                                        <= Join_ss_inst_ss_net_profit_bus_rdat_ready;
  Join_ss_inst_ss_store_sk_bus_rreq_ready                                                             <= RDAW64DW512LW8BS1BM16_inst_bsv_rreq_ready(3);
  Join_ss_inst_ss_store_sk_bus_rdat_valid                                                             <= RDAW64DW512LW8BS1BM16_inst_bsv_rdat_valid(3);
  Join_ss_inst_ss_store_sk_bus_rdat_last                                                              <= RDAW64DW512LW8BS1BM16_inst_bsv_rdat_last(3);
  Join_ss_inst_ss_store_sk_bus_rdat_data                                                              <= RDAW64DW512LW8BS1BM16_inst_bsv_rdat_data(BUS_DATA_WIDTH*3+BUS_DATA_WIDTH-1 downto BUS_DATA_WIDTH*3);
  Join_ss_inst_ss_sold_date_sk_bus_rreq_ready                                                         <= RDAW64DW512LW8BS1BM16_inst_bsv_rreq_ready(0);
  Join_ss_inst_ss_sold_date_sk_bus_rdat_valid                                                         <= RDAW64DW512LW8BS1BM16_inst_bsv_rdat_valid(0);
  Join_ss_inst_ss_sold_date_sk_bus_rdat_last                                                          <= RDAW64DW512LW8BS1BM16_inst_bsv_rdat_last(0);
  Join_ss_inst_ss_sold_date_sk_bus_rdat_data                                                          <= RDAW64DW512LW8BS1BM16_inst_bsv_rdat_data(BUS_DATA_WIDTH-1 downto 0);
  Join_ss_inst_ss_sales_price_bus_rreq_ready                                                          <= RDAW64DW512LW8BS1BM16_inst_bsv_rreq_ready(5);
  Join_ss_inst_ss_sales_price_bus_rdat_valid                                                          <= RDAW64DW512LW8BS1BM16_inst_bsv_rdat_valid(5);
  Join_ss_inst_ss_sales_price_bus_rdat_last                                                           <= RDAW64DW512LW8BS1BM16_inst_bsv_rdat_last(5);
  Join_ss_inst_ss_sales_price_bus_rdat_data                                                           <= RDAW64DW512LW8BS1BM16_inst_bsv_rdat_data(BUS_DATA_WIDTH*5+BUS_DATA_WIDTH-1 downto BUS_DATA_WIDTH*5);
  Join_ss_inst_ss_quantity_bus_rreq_ready                                                             <= RDAW64DW512LW8BS1BM16_inst_bsv_rreq_ready(4);
  Join_ss_inst_ss_quantity_bus_rdat_valid                                                             <= RDAW64DW512LW8BS1BM16_inst_bsv_rdat_valid(4);
  Join_ss_inst_ss_quantity_bus_rdat_last                                                              <= RDAW64DW512LW8BS1BM16_inst_bsv_rdat_last(4);
  Join_ss_inst_ss_quantity_bus_rdat_data                                                              <= RDAW64DW512LW8BS1BM16_inst_bsv_rdat_data(BUS_DATA_WIDTH*4+BUS_DATA_WIDTH-1 downto BUS_DATA_WIDTH*4);
  Join_ss_inst_ss_net_profit_bus_rreq_ready                                                           <= RDAW64DW512LW8BS1BM16_inst_bsv_rreq_ready(6);
  Join_ss_inst_ss_net_profit_bus_rdat_valid                                                           <= RDAW64DW512LW8BS1BM16_inst_bsv_rdat_valid(6);
  Join_ss_inst_ss_net_profit_bus_rdat_last                                                            <= RDAW64DW512LW8BS1BM16_inst_bsv_rdat_last(6);
  Join_ss_inst_ss_net_profit_bus_rdat_data                                                            <= RDAW64DW512LW8BS1BM16_inst_bsv_rdat_data(BUS_DATA_WIDTH*6+BUS_DATA_WIDTH-1 downto BUS_DATA_WIDTH*6);
  Join_ss_inst_ss_cdemo_sk_bus_rreq_ready                                                             <= RDAW64DW512LW8BS1BM16_inst_bsv_rreq_ready(1);
  Join_ss_inst_ss_cdemo_sk_bus_rdat_valid                                                             <= RDAW64DW512LW8BS1BM16_inst_bsv_rdat_valid(1);
  Join_ss_inst_ss_cdemo_sk_bus_rdat_last                                                              <= RDAW64DW512LW8BS1BM16_inst_bsv_rdat_last(1);
  Join_ss_inst_ss_cdemo_sk_bus_rdat_data                                                              <= RDAW64DW512LW8BS1BM16_inst_bsv_rdat_data(BUS_DATA_WIDTH+BUS_DATA_WIDTH-1 downto BUS_DATA_WIDTH);
  Join_ss_inst_ss_addr_sk_bus_rreq_ready                                                              <= RDAW64DW512LW8BS1BM16_inst_bsv_rreq_ready(2);
  Join_ss_inst_ss_addr_sk_bus_rdat_valid                                                              <= RDAW64DW512LW8BS1BM16_inst_bsv_rdat_valid(2);
  Join_ss_inst_ss_addr_sk_bus_rdat_last                                                               <= RDAW64DW512LW8BS1BM16_inst_bsv_rdat_last(2);
  Join_ss_inst_ss_addr_sk_bus_rdat_data                                                               <= RDAW64DW512LW8BS1BM16_inst_bsv_rdat_data(BUS_DATA_WIDTH*2+BUS_DATA_WIDTH-1 downto BUS_DATA_WIDTH*2);

end architecture;
