-- Copyright 2018-2019 Delft University of Technology
--
-- Licensed under the Apache License, Version 2.0 (the "License");
-- you may not use this file except in compliance with the License.
-- You may obtain a copy of the License at
--
--     http://www.apache.org/licenses/LICENSE-2.0
--
-- Unless required by applicable law or agreed to in writing, software
-- distributed under the License is distributed on an "AS IS" BASIS,
-- WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
-- See the License for the specific language governing permissions and
-- limitations under the License.
--
-- This file was generated by Fletchgen. Modify this file at your own risk.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity Join is
  generic (
    INDEX_WIDTH : integer := 32;
    TAG_WIDTH   : integer := 1
  );
  port (
    kcd_clk                      : in  std_logic;
    kcd_reset                    : in  std_logic;
    ss_sold_date_sk_valid        : in  std_logic;
    ss_sold_date_sk_ready        : out std_logic;
    ss_sold_date_sk_dvalid       : in  std_logic;
    ss_sold_date_sk_last         : in  std_logic;
    ss_sold_date_sk              : in  std_logic_vector(63 downto 0);
    ss_cdemo_sk_valid            : in  std_logic;
    ss_cdemo_sk_ready            : out std_logic;
    ss_cdemo_sk_dvalid           : in  std_logic;
    ss_cdemo_sk_last             : in  std_logic;
    ss_cdemo_sk                  : in  std_logic_vector(63 downto 0);
    ss_addr_sk_valid             : in  std_logic;
    ss_addr_sk_ready             : out std_logic;
    ss_addr_sk_dvalid            : in  std_logic;
    ss_addr_sk_last              : in  std_logic;
    ss_addr_sk                   : in  std_logic_vector(63 downto 0);
    ss_store_sk_valid            : in  std_logic;
    ss_store_sk_ready            : out std_logic;
    ss_store_sk_dvalid           : in  std_logic;
    ss_store_sk_last             : in  std_logic;
    ss_store_sk                  : in  std_logic_vector(63 downto 0);
    ss_quantity_valid            : in  std_logic;
    ss_quantity_ready            : out std_logic;
    ss_quantity_dvalid           : in  std_logic;
    ss_quantity_last             : in  std_logic;
    ss_quantity                  : in  std_logic_vector(63 downto 0);
    ss_sales_price_valid         : in  std_logic;
    ss_sales_price_ready         : out std_logic;
    ss_sales_price_dvalid        : in  std_logic;
    ss_sales_price_last          : in  std_logic;
    ss_sales_price               : in  std_logic_vector(63 downto 0);
    ss_net_profit_valid          : in  std_logic;
    ss_net_profit_ready          : out std_logic;
    ss_net_profit_dvalid         : in  std_logic;
    ss_net_profit_last           : in  std_logic;
    ss_net_profit                : in  std_logic_vector(63 downto 0);
    ss_sold_date_sk_unl_valid    : in  std_logic;
    ss_sold_date_sk_unl_ready    : out std_logic;
    ss_sold_date_sk_unl_tag      : in  std_logic_vector(TAG_WIDTH-1 downto 0);
    ss_cdemo_sk_unl_valid        : in  std_logic;
    ss_cdemo_sk_unl_ready        : out std_logic;
    ss_cdemo_sk_unl_tag          : in  std_logic_vector(TAG_WIDTH-1 downto 0);
    ss_addr_sk_unl_valid         : in  std_logic;
    ss_addr_sk_unl_ready         : out std_logic;
    ss_addr_sk_unl_tag           : in  std_logic_vector(TAG_WIDTH-1 downto 0);
    ss_store_sk_unl_valid        : in  std_logic;
    ss_store_sk_unl_ready        : out std_logic;
    ss_store_sk_unl_tag          : in  std_logic_vector(TAG_WIDTH-1 downto 0);
    ss_quantity_unl_valid        : in  std_logic;
    ss_quantity_unl_ready        : out std_logic;
    ss_quantity_unl_tag          : in  std_logic_vector(TAG_WIDTH-1 downto 0);
    ss_sales_price_unl_valid     : in  std_logic;
    ss_sales_price_unl_ready     : out std_logic;
    ss_sales_price_unl_tag       : in  std_logic_vector(TAG_WIDTH-1 downto 0);
    ss_net_profit_unl_valid      : in  std_logic;
    ss_net_profit_unl_ready      : out std_logic;
    ss_net_profit_unl_tag        : in  std_logic_vector(TAG_WIDTH-1 downto 0);
    ss_sold_date_sk_cmd_valid    : out std_logic;
    ss_sold_date_sk_cmd_ready    : in  std_logic;
    ss_sold_date_sk_cmd_firstIdx : out std_logic_vector(INDEX_WIDTH-1 downto 0);
    ss_sold_date_sk_cmd_lastIdx  : out std_logic_vector(INDEX_WIDTH-1 downto 0);
    ss_sold_date_sk_cmd_tag      : out std_logic_vector(TAG_WIDTH-1 downto 0);
    ss_cdemo_sk_cmd_valid        : out std_logic;
    ss_cdemo_sk_cmd_ready        : in  std_logic;
    ss_cdemo_sk_cmd_firstIdx     : out std_logic_vector(INDEX_WIDTH-1 downto 0);
    ss_cdemo_sk_cmd_lastIdx      : out std_logic_vector(INDEX_WIDTH-1 downto 0);
    ss_cdemo_sk_cmd_tag          : out std_logic_vector(TAG_WIDTH-1 downto 0);
    ss_addr_sk_cmd_valid         : out std_logic;
    ss_addr_sk_cmd_ready         : in  std_logic;
    ss_addr_sk_cmd_firstIdx      : out std_logic_vector(INDEX_WIDTH-1 downto 0);
    ss_addr_sk_cmd_lastIdx       : out std_logic_vector(INDEX_WIDTH-1 downto 0);
    ss_addr_sk_cmd_tag           : out std_logic_vector(TAG_WIDTH-1 downto 0);
    ss_store_sk_cmd_valid        : out std_logic;
    ss_store_sk_cmd_ready        : in  std_logic;
    ss_store_sk_cmd_firstIdx     : out std_logic_vector(INDEX_WIDTH-1 downto 0);
    ss_store_sk_cmd_lastIdx      : out std_logic_vector(INDEX_WIDTH-1 downto 0);
    ss_store_sk_cmd_tag          : out std_logic_vector(TAG_WIDTH-1 downto 0);
    ss_quantity_cmd_valid        : out std_logic;
    ss_quantity_cmd_ready        : in  std_logic;
    ss_quantity_cmd_firstIdx     : out std_logic_vector(INDEX_WIDTH-1 downto 0);
    ss_quantity_cmd_lastIdx      : out std_logic_vector(INDEX_WIDTH-1 downto 0);
    ss_quantity_cmd_tag          : out std_logic_vector(TAG_WIDTH-1 downto 0);
    ss_sales_price_cmd_valid     : out std_logic;
    ss_sales_price_cmd_ready     : in  std_logic;
    ss_sales_price_cmd_firstIdx  : out std_logic_vector(INDEX_WIDTH-1 downto 0);
    ss_sales_price_cmd_lastIdx   : out std_logic_vector(INDEX_WIDTH-1 downto 0);
    ss_sales_price_cmd_tag       : out std_logic_vector(TAG_WIDTH-1 downto 0);
    ss_net_profit_cmd_valid      : out std_logic;
    ss_net_profit_cmd_ready      : in  std_logic;
    ss_net_profit_cmd_firstIdx   : out std_logic_vector(INDEX_WIDTH-1 downto 0);
    ss_net_profit_cmd_lastIdx    : out std_logic_vector(INDEX_WIDTH-1 downto 0);
    ss_net_profit_cmd_tag        : out std_logic_vector(TAG_WIDTH-1 downto 0);
    start                        : in  std_logic;
    stop                         : in  std_logic;
    reset                        : in  std_logic;
    idle                         : out std_logic;
    busy                         : out std_logic;
    done                         : out std_logic;
    result                       : out std_logic_vector(63 downto 0);
    ss_firstidx                  : in  std_logic_vector(31 downto 0);
    ss_lastidx                   : in  std_logic_vector(31 downto 0)
  );
end entity;

architecture Implementation of Join is
begin
end architecture;
